* NGSPICE file created from TOP.ext - technology: gf180mcuD

.subckt TOP VDD VCTRL OUT VCNB VCNS VSS
X0 VDD.t17 a_n8471_219.t5 a_3149_2840 VDD.t16 pfet_03v3 ad=0.585p pd=3.1u as=0.585p ps=3.1u w=0.9u l=0.33u
X1 VSS.t18 a_n4208_n141.t3 a_n671_n1138 VSS.t0 nfet_03v3 ad=0.2646p pd=2.1u as=0.2646p ps=2.1u w=0.42u l=0.33u
X2 OUT.t1 a_11009_2840 a_14657_n1138 VSS.t15 nfet_03v3 ad=0.5124p pd=2.9u as=0.5124p ps=2.9u w=0.84u l=0.33u
X3 a_7177_2840 a_3345_2840 a_6981_2840 VDD.t18 pfet_03v3 ad=1.17p pd=4.9u as=1.17p ps=4.9u w=1.8u l=0.33u
X4 VSS.t4 VCNS.t0 a_n8659_n1230 VSS.t3 nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.33u
X5 VSS.t6 a_16431_6193 VSS.t5 ppolyf_u r_width=0.8u r_length=0.13m
X6 a_n8471_219.t0 VCNB.t0 a_n8659_n1230 VSS.t23 nfet_03v3 ad=0.52p pd=2.52u as=1.22p ps=5.22u w=2u l=0.33u
X7 VDD.t15 a_n8471_219.t6 a_18477_2840 VDD.t14 pfet_03v3 ad=0.585p pd=3.1u as=0.585p ps=3.1u w=0.9u l=0.33u
X8 VSS.t24 VCNS.t1 a_n8659_n1230 VSS.t23 nfet_03v3 ad=0.52p pd=2.52u as=1.22p ps=5.22u w=2u l=0.33u
X9 VDD.t13 a_n8471_219.t1 a_n8471_219.t2 VDD.t12 pfet_03v3 ad=0.585p pd=3.1u as=0.585p ps=3.1u w=0.9u l=0.33u
X10 VDD.t11 a_n8471_219.t7 a_n683_2840 VDD.t10 pfet_03v3 ad=0.585p pd=3.1u as=0.585p ps=3.1u w=0.9u l=0.33u
X11 a_11009_2840 a_7177_2840 a_10813_2840 VDD.t21 pfet_03v3 ad=1.17p pd=4.9u as=1.17p ps=4.9u w=1.8u l=0.33u
X12 a_3345_2840 a_n487_2840 a_3149_2840 VDD.t20 pfet_03v3 ad=1.17p pd=4.9u as=1.17p ps=4.9u w=1.8u l=0.33u
X13 a_n4208_n141.t0 a_n8471_219.t8 VDD.t9 VDD.t8 pfet_03v3 ad=0.585p pd=3.1u as=0.585p ps=3.1u w=0.9u l=0.33u
X14 a_n487_2840 OUT.t2 a_n671_n1138 VSS.t0 nfet_03v3 ad=0.5124p pd=2.9u as=0.5124p ps=2.9u w=0.84u l=0.33u
X15 a_7177_2840 a_3345_2840 a_6993_n1138 VSS.t9 nfet_03v3 ad=0.5124p pd=2.9u as=0.5124p ps=2.9u w=0.84u l=0.33u
X16 a_n8471_219.t4 VCTRL.t0 a_n9701_6193 VSS.t22 nfet_03v3 ad=0.488p pd=2.82u as=0.488p ps=2.82u w=0.8u l=0.33u
X17 a_18673_2840 OUT.t3 a_18477_2840 VDD.t0 pfet_03v3 ad=1.17p pd=4.9u as=1.17p ps=4.9u w=1.8u l=0.33u
X18 a_18673_2840 OUT.t4 a_18489_n1138 VSS.t2 nfet_03v3 ad=0.5124p pd=2.9u as=0.5124p ps=2.9u w=0.84u l=0.33u
X19 VSS.t17 a_n4208_n141.t4 a_18489_n1138 VSS.t2 nfet_03v3 ad=0.2646p pd=2.1u as=0.2646p ps=2.1u w=0.42u l=0.33u
X20 a_n487_2840 OUT.t5 a_n683_2840 VDD.t1 pfet_03v3 ad=1.17p pd=4.9u as=1.17p ps=4.9u w=1.8u l=0.33u
X21 a_n8659_n1230 VCNS.t2 VSS.t21 VSS.t1 nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.33u
X22 VDD.t7 a_n8471_219.t9 a_14645_2840 VDD.t6 pfet_03v3 ad=0.585p pd=3.1u as=0.585p ps=3.1u w=0.9u l=0.33u
X23 VSS.t16 a_n4208_n141.t5 a_14657_n1138 VSS.t15 nfet_03v3 ad=0.2646p pd=2.1u as=0.2646p ps=2.1u w=0.42u l=0.33u
X24 VSS.t14 a_n4208_n141.t6 a_3161_n1138 VSS.t13 nfet_03v3 ad=0.2646p pd=2.1u as=0.2646p ps=2.1u w=0.42u l=0.33u
X25 VDD.t5 a_n8471_219.t10 a_6981_2840 VDD.t4 pfet_03v3 ad=0.585p pd=3.1u as=0.585p ps=3.1u w=0.9u l=0.33u
X26 a_n8471_219.t3 VCNB.t1 a_n8659_n1230 VSS.t3 nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.33u
X27 a_n4208_n141.t2 a_n4208_n141.t1 VSS.t12 VSS.t11 nfet_03v3 ad=0.2646p pd=2.1u as=0.2646p ps=2.1u w=0.42u l=0.33u
X28 a_11009_2840 a_7177_2840 a_10825_n1138 VSS.t7 nfet_03v3 ad=0.5124p pd=2.9u as=0.5124p ps=2.9u w=0.84u l=0.33u
X29 VSS.t10 a_n4208_n141.t7 a_6993_n1138 VSS.t9 nfet_03v3 ad=0.2646p pd=2.1u as=0.2646p ps=2.1u w=0.42u l=0.33u
X30 a_n8659_n1230 VCNB.t2 a_n8471_219.t3 VSS.t19 nfet_03v3 ad=1.22p pd=5.22u as=0.52p ps=2.52u w=2u l=0.33u
X31 a_n8659_n1230 VCNS.t3 VSS.t20 VSS.t19 nfet_03v3 ad=1.22p pd=5.22u as=0.52p ps=2.52u w=2u l=0.33u
X32 a_3345_2840 a_n487_2840 a_3161_n1138 VSS.t13 nfet_03v3 ad=0.5124p pd=2.9u as=0.5124p ps=2.9u w=0.84u l=0.33u
X33 VSS.t8 a_n4208_n141.t8 a_10825_n1138 VSS.t7 nfet_03v3 ad=0.2646p pd=2.1u as=0.2646p ps=2.1u w=0.42u l=0.33u
X34 a_n9701_6193 a_16431_6193 VSS.t5 ppolyf_u r_width=0.8u r_length=0.13m
X35 VDD.t3 a_n8471_219.t11 a_10813_2840 VDD.t2 pfet_03v3 ad=0.585p pd=3.1u as=0.585p ps=3.1u w=0.9u l=0.33u
X36 a_n8659_n1230 VCNB.t3 a_n8471_219.t0 VSS.t1 nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.33u
X37 OUT.t0 a_11009_2840 a_14645_2840 VDD.t19 pfet_03v3 ad=1.17p pd=4.9u as=1.17p ps=4.9u w=1.8u l=0.33u
R0 a_n8471_219.n1 a_n8471_219.t6 31.1854
R1 a_n8471_219.n0 a_n8471_219.t8 30.4809
R2 a_n8471_219.n0 a_n8471_219.t7 29.7468
R3 a_n8471_219.n0 a_n8471_219.t5 29.7468
R4 a_n8471_219.n2 a_n8471_219.t10 29.7468
R5 a_n8471_219.n2 a_n8471_219.t11 29.7468
R6 a_n8471_219.n1 a_n8471_219.t9 29.7468
R7 a_n8471_219.n3 a_n8471_219.t1 28.2414
R8 a_n8471_219.n0 a_n8471_219.t4 11.7439
R9 a_n8471_219.n3 a_n8471_219.t2 8.52921
R10 a_n8471_219.t0 a_n8471_219.n4 4.56638
R11 a_n8471_219.n4 a_n8471_219.t3 4.38259
R12 a_n8471_219.n4 a_n8471_219.n0 3.5234
R13 a_n8471_219.n0 a_n8471_219.n2 2.8778
R14 a_n8471_219.n2 a_n8471_219.n1 2.8778
R15 a_n8471_219.n0 a_n8471_219.n3 2.4541
R16 VDD.n2 VDD.t14 589.355
R17 VDD.n8 VDD.t6 589.355
R18 VDD.n15 VDD.t2 589.355
R19 VDD.n22 VDD.t4 589.355
R20 VDD.n29 VDD.t16 589.355
R21 VDD.n36 VDD.t10 589.355
R22 VDD.n42 VDD.t12 589.355
R23 VDD.n41 VDD.t8 589.355
R24 VDD.n3 VDD.t0 419.211
R25 VDD.n9 VDD.t19 419.211
R26 VDD.n16 VDD.t21 419.211
R27 VDD.n23 VDD.t18 419.211
R28 VDD.n30 VDD.t20 419.211
R29 VDD.n37 VDD.t1 419.211
R30 VDD.n42 VDD.t13 8.52192
R31 VDD.n41 VDD.t9 8.52192
R32 VDD.n2 VDD.t15 8.46717
R33 VDD.n8 VDD.t7 8.46717
R34 VDD.n15 VDD.t3 8.46717
R35 VDD.n22 VDD.t5 8.46717
R36 VDD.n29 VDD.t17 8.46717
R37 VDD.n36 VDD.t11 8.46717
R38 VDD.n4 VDD.n1 4.5005
R39 VDD.n1 VDD.n0 4.5005
R40 VDD.n4 VDD.n3 4.5005
R41 VDD.n3 VDD.n0 4.5005
R42 VDD.n10 VDD.n7 4.5005
R43 VDD.n7 VDD.n6 4.5005
R44 VDD.n10 VDD.n9 4.5005
R45 VDD.n9 VDD.n6 4.5005
R46 VDD.n17 VDD.n14 4.5005
R47 VDD.n14 VDD.n13 4.5005
R48 VDD.n17 VDD.n16 4.5005
R49 VDD.n16 VDD.n13 4.5005
R50 VDD.n24 VDD.n21 4.5005
R51 VDD.n21 VDD.n20 4.5005
R52 VDD.n24 VDD.n23 4.5005
R53 VDD.n23 VDD.n20 4.5005
R54 VDD.n31 VDD.n28 4.5005
R55 VDD.n28 VDD.n27 4.5005
R56 VDD.n31 VDD.n30 4.5005
R57 VDD.n30 VDD.n27 4.5005
R58 VDD.n38 VDD.n35 4.5005
R59 VDD.n35 VDD.n34 4.5005
R60 VDD.n38 VDD.n37 4.5005
R61 VDD.n37 VDD.n34 4.5005
R62 VDD.n44 VDD.n43 4.06871
R63 VDD VDD.n5 3.40475
R64 VDD.n12 VDD.n11 2.70462
R65 VDD.n19 VDD.n18 2.70462
R66 VDD.n26 VDD.n25 2.70462
R67 VDD.n33 VDD.n32 2.70462
R68 VDD.n40 VDD.n39 2.70462
R69 VDD VDD.n44 0.777875
R70 VDD.n12 VDD 0.737375
R71 VDD.n19 VDD 0.7265
R72 VDD.n26 VDD 0.7265
R73 VDD.n33 VDD 0.7265
R74 VDD.n40 VDD 0.7265
R75 VDD.n44 VDD 0.7265
R76 VDD VDD.n12 0.7115
R77 VDD VDD.n19 0.7115
R78 VDD VDD.n26 0.7115
R79 VDD VDD.n33 0.7115
R80 VDD VDD.n40 0.7115
R81 VDD.n43 VDD.n42 0.181952
R82 VDD.n43 VDD.n41 0.146702
R83 VDD.n5 VDD.n4 0.024117
R84 VDD.n11 VDD.n10 0.024117
R85 VDD.n18 VDD.n17 0.024117
R86 VDD.n25 VDD.n24 0.024117
R87 VDD.n32 VDD.n31 0.024117
R88 VDD.n39 VDD.n38 0.024117
R89 VDD.n5 VDD.n0 0.0237979
R90 VDD.n11 VDD.n6 0.0237979
R91 VDD.n18 VDD.n13 0.0237979
R92 VDD.n25 VDD.n20 0.0237979
R93 VDD.n32 VDD.n27 0.0237979
R94 VDD.n39 VDD.n34 0.0237979
R95 VDD.n2 VDD.n1 0.020375
R96 VDD.n3 VDD.n2 0.020375
R97 VDD.n8 VDD.n7 0.020375
R98 VDD.n9 VDD.n8 0.020375
R99 VDD.n15 VDD.n14 0.020375
R100 VDD.n16 VDD.n15 0.020375
R101 VDD.n22 VDD.n21 0.020375
R102 VDD.n23 VDD.n22 0.020375
R103 VDD.n29 VDD.n28 0.020375
R104 VDD.n30 VDD.n29 0.020375
R105 VDD.n36 VDD.n35 0.020375
R106 VDD.n37 VDD.n36 0.020375
R107 a_n4208_n141.n2 a_n4208_n141.t4 26.5147
R108 a_n4208_n141.n1 a_n4208_n141.t3 25.076
R109 a_n4208_n141.n1 a_n4208_n141.t6 25.076
R110 a_n4208_n141.n3 a_n4208_n141.t7 25.076
R111 a_n4208_n141.n3 a_n4208_n141.t8 25.076
R112 a_n4208_n141.n2 a_n4208_n141.t5 25.076
R113 a_n4208_n141.n0 a_n4208_n141.t1 23.009
R114 a_n4208_n141.n0 a_n4208_n141.t2 12.3005
R115 a_n4208_n141.t0 a_n4208_n141.n1 11.2556
R116 a_n4208_n141.n1 a_n4208_n141.n0 3.08843
R117 a_n4208_n141.n1 a_n4208_n141.n3 2.8778
R118 a_n4208_n141.n3 a_n4208_n141.n2 2.8778
R119 VSS.n1905 VSS.n1904 30440.7
R120 VSS.n1904 VSS.n1886 21018.6
R121 VSS.n1905 VSS.n234 17216.6
R122 VSS.n1886 VSS.n234 11887.6
R123 VSS.n207 VSS.t22 8334.77
R124 VSS.n1953 VSS.n1952 6332.65
R125 VSS.n2063 VSS.n2062 6053.81
R126 VSS.n1904 VSS.n235 5872.22
R127 VSS.n1904 VSS.n1903 4786.34
R128 VSS.n1820 VSS.n234 4237.55
R129 VSS.n142 VSS.n138 3851.03
R130 VSS.n1821 VSS.n234 3453.21
R131 VSS.n778 VSS.n197 2950.24
R132 VSS.n1045 VSS.n1044 2950.24
R133 VSS.n778 VSS.n318 2950.24
R134 VSS.n1629 VSS.n318 2950.24
R135 VSS.n1629 VSS.n259 2950.24
R136 VSS.n1774 VSS.n259 2950.24
R137 VSS.n2294 VSS.n2293 2713.07
R138 VSS.n206 VSS.n205 2388.26
R139 VSS.n2062 VSS.t5 2153.74
R140 VSS.n976 VSS.n197 1959.56
R141 VSS.n941 VSS.n197 1959.56
R142 VSS.n1737 VSS.n197 1959.56
R143 VSS.n906 VSS.n197 1959.56
R144 VSS.n1654 VSS.n197 1959.56
R145 VSS.n2062 VSS.n196 1873.92
R146 VSS.n2212 VSS.n142 1727.25
R147 VSS.n746 VSS.n740 781.367
R148 VSS.n206 VSS.n142 659.034
R149 VSS.t5 VSS.n2061 623.524
R150 VSS.n2061 VSS.n199 621.324
R151 VSS.n2293 VSS.n45 551.149
R152 VSS.n2271 VSS.n45 504.923
R153 VSS.n2263 VSS.n2262 487.846
R154 VSS.n1549 VSS.n1548 487.846
R155 VSS.n453 VSS.n452 487.846
R156 VSS.n1362 VSS.n502 487.846
R157 VSS.n1234 VSS.n556 487.846
R158 VSS.n1106 VSS.n610 487.846
R159 VSS.n207 VSS.n196 475.474
R160 VSS.n716 VSS.n197 475.276
R161 VSS.n826 VSS.n197 475.276
R162 VSS.n1646 VSS.n197 475.276
R163 VSS.n1729 VSS.n197 475.276
R164 VSS.n1549 VSS.n359 461.786
R165 VSS.n452 VSS.n433 461.786
R166 VSS.n1363 VSS.n1362 461.786
R167 VSS.n1235 VSS.n1234 461.786
R168 VSS.n1107 VSS.n1106 461.786
R169 VSS.n198 VSS.n197 429.887
R170 VSS.n1555 VSS.n359 425.95
R171 VSS.n1556 VSS.n1555 425.95
R172 VSS.n1557 VSS.n1556 425.95
R173 VSS.n1557 VSS.n355 425.95
R174 VSS.n1563 VSS.n355 425.95
R175 VSS.n1564 VSS.n1563 425.95
R176 VSS.n1565 VSS.n1564 425.95
R177 VSS.n1565 VSS.n351 425.95
R178 VSS.n1571 VSS.n8 425.95
R179 VSS.n2356 VSS.n8 425.95
R180 VSS.n2254 VSS.n9 425.95
R181 VSS.n2255 VSS.n2254 425.95
R182 VSS.n2255 VSS.n2251 425.95
R183 VSS.n2261 VSS.n2251 425.95
R184 VSS.n2262 VSS.n2261 425.95
R185 VSS.n1516 VSS.n433 425.95
R186 VSS.n1517 VSS.n1516 425.95
R187 VSS.n1518 VSS.n1517 425.95
R188 VSS.n1518 VSS.n429 425.95
R189 VSS.n1524 VSS.n429 425.95
R190 VSS.n1525 VSS.n1524 425.95
R191 VSS.n1527 VSS.n1525 425.95
R192 VSS.n1527 VSS.n1526 425.95
R193 VSS.n1534 VSS.n1533 425.95
R194 VSS.n1535 VSS.n1534 425.95
R195 VSS.n1540 VSS.n1539 425.95
R196 VSS.n1541 VSS.n1540 425.95
R197 VSS.n1541 VSS.n363 425.95
R198 VSS.n1547 VSS.n363 425.95
R199 VSS.n1548 VSS.n1547 425.95
R200 VSS.n1384 VSS.n1363 425.95
R201 VSS.n1384 VSS.n1383 425.95
R202 VSS.n1383 VSS.n1382 425.95
R203 VSS.n1382 VSS.n1364 425.95
R204 VSS.n1376 VSS.n1364 425.95
R205 VSS.n1376 VSS.n1375 425.95
R206 VSS.n1375 VSS.n1374 425.95
R207 VSS.n1374 VSS.n487 425.95
R208 VSS.n488 VSS.n444 425.95
R209 VSS.n1509 VSS.n444 425.95
R210 VSS.n462 VSS.n461 425.95
R211 VSS.n461 VSS.n445 425.95
R212 VSS.n449 VSS.n445 425.95
R213 VSS.n454 VSS.n449 425.95
R214 VSS.n454 VSS.n453 425.95
R215 VSS.n1256 VSS.n1235 425.95
R216 VSS.n1256 VSS.n1255 425.95
R217 VSS.n1255 VSS.n1254 425.95
R218 VSS.n1254 VSS.n1236 425.95
R219 VSS.n1248 VSS.n1236 425.95
R220 VSS.n1248 VSS.n1247 425.95
R221 VSS.n1247 VSS.n1246 425.95
R222 VSS.n1246 VSS.n540 425.95
R223 VSS.n541 VSS.n514 425.95
R224 VSS.n1348 VSS.n514 425.95
R225 VSS.n515 VSS.n506 425.95
R226 VSS.n1354 VSS.n506 425.95
R227 VSS.n1355 VSS.n1354 425.95
R228 VSS.n1356 VSS.n1355 425.95
R229 VSS.n1356 VSS.n502 425.95
R230 VSS.n1128 VSS.n1107 425.95
R231 VSS.n1128 VSS.n1127 425.95
R232 VSS.n1127 VSS.n1126 425.95
R233 VSS.n1126 VSS.n1108 425.95
R234 VSS.n1120 VSS.n1108 425.95
R235 VSS.n1120 VSS.n1119 425.95
R236 VSS.n1119 VSS.n1118 425.95
R237 VSS.n1118 VSS.n594 425.95
R238 VSS.n595 VSS.n568 425.95
R239 VSS.n1220 VSS.n568 425.95
R240 VSS.n569 VSS.n560 425.95
R241 VSS.n1226 VSS.n560 425.95
R242 VSS.n1227 VSS.n1226 425.95
R243 VSS.n1228 VSS.n1227 425.95
R244 VSS.n1228 VSS.n556 425.95
R245 VSS.n1092 VSS.n614 425.95
R246 VSS.n1098 VSS.n614 425.95
R247 VSS.n1099 VSS.n1098 425.95
R248 VSS.n1100 VSS.n1099 425.95
R249 VSS.n1100 VSS.n610 425.95
R250 VSS.n1953 VSS.n198 350.44
R251 VSS.n2029 VSS.n2028 302.466
R252 VSS.n2028 VSS.n2027 302.466
R253 VSS.n2027 VSS.n1986 302.466
R254 VSS.n2021 VSS.n1986 302.466
R255 VSS.n2021 VSS.n2020 302.466
R256 VSS.n2020 VSS.n2019 302.466
R257 VSS.n2019 VSS.n1991 302.466
R258 VSS.n2013 VSS.n1991 302.466
R259 VSS.n747 VSS.n746 278.373
R260 VSS.n747 VSS.n685 278.373
R261 VSS.n1758 VSS.n264 272.08
R262 VSS.n1764 VSS.n264 272.08
R263 VSS.n1765 VSS.n1764 272.08
R264 VSS.n1766 VSS.n1765 272.08
R265 VSS.n1766 VSS.n260 272.08
R266 VSS.n1772 VSS.n260 272.08
R267 VSS.n1773 VSS.n1772 272.08
R268 VSS.n1775 VSS.n255 272.08
R269 VSS.n1781 VSS.n255 272.08
R270 VSS.n1782 VSS.n1781 272.08
R271 VSS.n1783 VSS.n1782 272.08
R272 VSS.n1783 VSS.n251 272.08
R273 VSS.n1789 VSS.n251 272.08
R274 VSS.n1790 VSS.n1789 272.08
R275 VSS.n1791 VSS.n1790 272.08
R276 VSS.n1838 VSS.n1837 272.08
R277 VSS.n1839 VSS.n1838 272.08
R278 VSS.n1839 VSS.n243 272.08
R279 VSS.n1845 VSS.n243 272.08
R280 VSS.n1846 VSS.n1845 272.08
R281 VSS.n1848 VSS.n236 272.08
R282 VSS.n1885 VSS.n237 272.08
R283 VSS.n1879 VSS.n237 272.08
R284 VSS.n1879 VSS.n1878 272.08
R285 VSS.n1878 VSS.n1877 272.08
R286 VSS.n1877 VSS.n1854 272.08
R287 VSS.n1871 VSS.n1854 272.08
R288 VSS.n1871 VSS.n1870 272.08
R289 VSS.n1870 VSS.n1869 272.08
R290 VSS.n1869 VSS.n1858 272.08
R291 VSS.n1863 VSS.n1858 272.08
R292 VSS.n1863 VSS.n1862 272.08
R293 VSS.n1862 VSS.n46 272.08
R294 VSS.n2355 VSS.n9 264.089
R295 VSS.n1539 VSS.n367 264.089
R296 VSS.n1508 VSS.n462 264.089
R297 VSS.n1347 VSS.n515 264.089
R298 VSS.n1219 VSS.n569 264.089
R299 VSS.n1847 VSS.n1846 263.918
R300 VSS.n1044 VSS.n685 250.536
R301 VSS.n739 VSS.n738 242.81
R302 VSS.n738 VSS.n724 242.81
R303 VSS.n732 VSS.n724 242.81
R304 VSS.n732 VSS.n731 242.81
R305 VSS.n731 VSS.n730 242.81
R306 VSS.n730 VSS.n684 242.81
R307 VSS.n1046 VSS.n684 242.81
R308 VSS.n1052 VSS.n680 242.81
R309 VSS.n1053 VSS.n1052 242.81
R310 VSS.n1055 VSS.n1053 242.81
R311 VSS.n1055 VSS.n1054 242.81
R312 VSS.n2293 VSS.n2292 235.351
R313 VSS.n1572 VSS.n1571 230.013
R314 VSS.n2356 VSS.n2355 230.013
R315 VSS.n1533 VSS.n425 230.013
R316 VSS.n1535 VSS.n367 230.013
R317 VSS.n1405 VSS.n488 230.013
R318 VSS.n1509 VSS.n1508 230.013
R319 VSS.n1277 VSS.n541 230.013
R320 VSS.n1348 VSS.n1347 230.013
R321 VSS.n1149 VSS.n595 230.013
R322 VSS.n1220 VSS.n1219 230.013
R323 VSS.n2068 VSS.n192 225.93
R324 VSS.n2069 VSS.n2068 225.93
R325 VSS.n2070 VSS.n2069 225.93
R326 VSS.n2070 VSS.n188 225.93
R327 VSS.n2076 VSS.n188 225.93
R328 VSS.n2081 VSS.n2079 225.93
R329 VSS.n2081 VSS.n2080 225.93
R330 VSS.n2061 VSS.n2060 216.263
R331 VSS.n811 VSS.n810 210.766
R332 VSS.n810 VSS.n809 210.766
R333 VSS.n809 VSS.n770 210.766
R334 VSS.n803 VSS.n770 210.766
R335 VSS.n803 VSS.n802 210.766
R336 VSS.n802 VSS.n801 210.766
R337 VSS.n801 VSS.n774 210.766
R338 VSS.n795 VSS.n794 210.766
R339 VSS.n794 VSS.n793 210.766
R340 VSS.n793 VSS.n779 210.766
R341 VSS.n787 VSS.n779 210.766
R342 VSS.n874 VSS.n873 210.766
R343 VSS.n873 VSS.n872 210.766
R344 VSS.n872 VSS.n834 210.766
R345 VSS.n866 VSS.n834 210.766
R346 VSS.n866 VSS.n865 210.766
R347 VSS.n865 VSS.n864 210.766
R348 VSS.n864 VSS.n838 210.766
R349 VSS.n858 VSS.n857 210.766
R350 VSS.n857 VSS.n856 210.766
R351 VSS.n856 VSS.n842 210.766
R352 VSS.n850 VSS.n842 210.766
R353 VSS.n1645 VSS.n306 210.766
R354 VSS.n1639 VSS.n306 210.766
R355 VSS.n1639 VSS.n1638 210.766
R356 VSS.n1638 VSS.n1637 210.766
R357 VSS.n1637 VSS.n314 210.766
R358 VSS.n1631 VSS.n314 210.766
R359 VSS.n1631 VSS.n1630 210.766
R360 VSS.n1628 VSS.n319 210.766
R361 VSS.n1622 VSS.n319 210.766
R362 VSS.n1622 VSS.n1621 210.766
R363 VSS.n1621 VSS.n1620 210.766
R364 VSS.n1728 VSS.n282 210.766
R365 VSS.n1722 VSS.n282 210.766
R366 VSS.n1722 VSS.n1721 210.766
R367 VSS.n1721 VSS.n1720 210.766
R368 VSS.n1720 VSS.n1688 210.766
R369 VSS.n1714 VSS.n1688 210.766
R370 VSS.n1714 VSS.n1713 210.766
R371 VSS.n1710 VSS.n1709 210.766
R372 VSS.n1709 VSS.n1708 210.766
R373 VSS.n1708 VSS.n1693 210.766
R374 VSS.n1702 VSS.n1693 210.766
R375 VSS.n2062 VSS.n192 208.986
R376 VSS.n1572 VSS.n351 195.938
R377 VSS.n1526 VSS.n425 195.938
R378 VSS.n1405 VSS.n487 195.938
R379 VSS.n1277 VSS.n540 195.938
R380 VSS.n1149 VSS.n594 195.938
R381 VSS.n1886 VSS.n236 195.899
R382 VSS.n218 VSS.n198 183.655
R383 VSS.n2263 VSS.n45 176.399
R384 VSS.n1775 VSS.n1774 168.69
R385 VSS.n2292 VSS.n47 168.69
R386 VSS.n1092 VSS.n1091 168.25
R387 VSS.n1837 VSS.n247 167.329
R388 VSS.n1084 VSS.n1070 157.006
R389 VSS.n1084 VSS.n1083 157.006
R390 VSS.n1083 VSS.n1082 157.006
R391 VSS.n1082 VSS.n1071 157.006
R392 VSS.n1076 VSS.n1071 157.006
R393 VSS.n1076 VSS.n1075 157.006
R394 VSS.n1075 VSS.n604 157.006
R395 VSS.n1139 VSS.n600 157.006
R396 VSS.n1140 VSS.n1139 157.006
R397 VSS.n1141 VSS.n1140 157.006
R398 VSS.n1141 VSS.n596 157.006
R399 VSS.n1148 VSS.n596 157.006
R400 VSS.n1151 VSS.n1150 157.006
R401 VSS.n1151 VSS.n577 157.006
R402 VSS.n1176 VSS.n1175 157.006
R403 VSS.n1175 VSS.n1174 157.006
R404 VSS.n1174 VSS.n1157 157.006
R405 VSS.n1168 VSS.n1157 157.006
R406 VSS.n1168 VSS.n1167 157.006
R407 VSS.n1167 VSS.n1166 157.006
R408 VSS.n1166 VSS.n1161 157.006
R409 VSS.n1161 VSS.n550 157.006
R410 VSS.n1267 VSS.n546 157.006
R411 VSS.n1268 VSS.n1267 157.006
R412 VSS.n1269 VSS.n1268 157.006
R413 VSS.n1269 VSS.n542 157.006
R414 VSS.n1276 VSS.n542 157.006
R415 VSS.n1279 VSS.n1278 157.006
R416 VSS.n1279 VSS.n523 157.006
R417 VSS.n1304 VSS.n1303 157.006
R418 VSS.n1303 VSS.n1302 157.006
R419 VSS.n1302 VSS.n1285 157.006
R420 VSS.n1296 VSS.n1285 157.006
R421 VSS.n1296 VSS.n1295 157.006
R422 VSS.n1295 VSS.n1294 157.006
R423 VSS.n1294 VSS.n1289 157.006
R424 VSS.n1289 VSS.n497 157.006
R425 VSS.n1395 VSS.n493 157.006
R426 VSS.n1396 VSS.n1395 157.006
R427 VSS.n1397 VSS.n1396 157.006
R428 VSS.n1397 VSS.n489 157.006
R429 VSS.n1404 VSS.n489 157.006
R430 VSS.n1407 VSS.n1406 157.006
R431 VSS.n1407 VSS.n470 157.006
R432 VSS.n1465 VSS.n1464 157.006
R433 VSS.n1464 VSS.n1463 157.006
R434 VSS.n1463 VSS.n1413 157.006
R435 VSS.n1457 VSS.n1413 157.006
R436 VSS.n1457 VSS.n1456 157.006
R437 VSS.n1456 VSS.n1455 157.006
R438 VSS.n1455 VSS.n1417 157.006
R439 VSS.n1449 VSS.n1417 157.006
R440 VSS.n1446 VSS.n1421 157.006
R441 VSS.n1440 VSS.n1421 157.006
R442 VSS.n1440 VSS.n1439 157.006
R443 VSS.n1439 VSS.n1438 157.006
R444 VSS.n1438 VSS.n1425 157.006
R445 VSS.n1432 VSS.n1431 157.006
R446 VSS.n1431 VSS.n1430 157.006
R447 VSS.n1607 VSS.n1606 157.006
R448 VSS.n1606 VSS.n1605 157.006
R449 VSS.n1605 VSS.n333 157.006
R450 VSS.n1599 VSS.n333 157.006
R451 VSS.n1599 VSS.n1598 157.006
R452 VSS.n1598 VSS.n1597 157.006
R453 VSS.n1597 VSS.n337 157.006
R454 VSS.n1591 VSS.n337 157.006
R455 VSS.n1588 VSS.n342 157.006
R456 VSS.n1582 VSS.n342 157.006
R457 VSS.n1582 VSS.n1581 157.006
R458 VSS.n1581 VSS.n1580 157.006
R459 VSS.n1580 VSS.n346 157.006
R460 VSS.n1574 VSS.n1573 157.006
R461 VSS.n1573 VSS.n17 157.006
R462 VSS.n2312 VSS.n2311 157.006
R463 VSS.n2311 VSS.n2310 157.006
R464 VSS.n2310 VSS.n35 157.006
R465 VSS.n2304 VSS.n35 157.006
R466 VSS.n2304 VSS.n2303 157.006
R467 VSS.n2303 VSS.n2302 157.006
R468 VSS.n2302 VSS.n39 157.006
R469 VSS.n2296 VSS.n39 157.006
R470 VSS.n1043 VSS.n686 152.905
R471 VSS.n1037 VSS.n686 152.905
R472 VSS.n1037 VSS.n1036 152.905
R473 VSS.n1036 VSS.n1035 152.905
R474 VSS.n1035 VSS.n692 152.905
R475 VSS.n1029 VSS.n692 152.905
R476 VSS.n1029 VSS.n1028 152.905
R477 VSS.n992 VSS.n991 152.905
R478 VSS.n991 VSS.n990 152.905
R479 VSS.n990 VSS.n704 152.905
R480 VSS.n984 VSS.n704 152.905
R481 VSS.n984 VSS.n983 152.905
R482 VSS.n983 VSS.n982 152.905
R483 VSS.n982 VSS.n709 152.905
R484 VSS.n1133 VSS.n1132 150.726
R485 VSS.n1261 VSS.n1260 150.726
R486 VSS.n1389 VSS.n1388 150.726
R487 VSS.n1448 VSS.n1447 150.726
R488 VSS.n1590 VSS.n1589 150.726
R489 VSS.n1045 VSS.n680 150.542
R490 VSS.n1054 VSS.n620 150.542
R491 VSS.n1758 VSS.n218 146.923
R492 VSS.n1847 VSS.n242 131.885
R493 VSS.n740 VSS.n739 131.118
R494 VSS.n795 VSS.n778 130.674
R495 VSS.n787 VSS.n533 130.674
R496 VSS.n858 VSS.n318 130.674
R497 VSS.n850 VSS.n480 130.674
R498 VSS.n1629 VSS.n1628 130.674
R499 VSS.n1620 VSS.n323 130.674
R500 VSS.n1710 VSS.n259 130.674
R501 VSS.n1702 VSS.n27 130.674
R502 VSS.n2060 VSS.n207 128.548
R503 VSS.n2013 VSS.n2012 120.987
R504 VSS.n2078 VSS.n2076 120.873
R505 VSS.n2090 VSS.n180 117.484
R506 VSS.n811 VSS.n716 113.814
R507 VSS.n874 VSS.n826 113.814
R508 VSS.n1646 VSS.n1645 113.814
R509 VSS.n1729 VSS.n1728 113.814
R510 VSS.t2 VSS.n600 107.549
R511 VSS.t15 VSS.n546 107.549
R512 VSS.t7 VSS.n493 107.549
R513 VSS.t9 VSS.n1446 107.549
R514 VSS.t13 VSS.n1588 107.549
R515 VSS.n242 VSS.t0 107.549
R516 VSS.n2079 VSS.n2078 105.058
R517 VSS.n1791 VSS.n247 104.751
R518 VSS.n1774 VSS.n1773 103.391
R519 VSS.n1091 VSS.n618 95.8393
R520 VSS.n1176 VSS.n587 95.7734
R521 VSS.n1304 VSS.n533 95.7734
R522 VSS.n1465 VSS.n480 95.7734
R523 VSS.n1607 VSS.n323 95.7734
R524 VSS.n2312 VSS.n27 95.7734
R525 VSS.n1150 VSS.n1149 94.2034
R526 VSS.n1278 VSS.n1277 94.2034
R527 VSS.n1406 VSS.n1405 94.2034
R528 VSS.n1432 VSS.n425 94.2034
R529 VSS.n1574 VSS.n1572 94.2034
R530 VSS.n1947 VSS.n229 93.8561
R531 VSS.n1914 VSS.n1913 93.8561
R532 VSS.n1941 VSS.n1940 93.8561
R533 VSS.n1922 VSS.n1915 93.8561
R534 VSS.n1934 VSS.n1923 93.8561
R535 VSS.n1933 VSS.n1924 93.8561
R536 VSS.n1927 VSS.n1926 93.8561
R537 VSS.n2237 VSS.n62 93.8561
R538 VSS.n2230 VSS.n2229 93.8561
R539 VSS.n2226 VSS.n127 93.8561
R540 VSS.n2225 VSS.n130 93.8561
R541 VSS.n135 VSS.n134 93.8561
R542 VSS.n2219 VSS.n2218 93.8561
R543 VSS.n1070 VSS.n620 92.6334
R544 VSS.n1046 VSS.n1045 92.268
R545 VSS.n2202 VSS.n2201 86.7903
R546 VSS.n2195 VSS.n158 86.7903
R547 VSS.n2194 VSS.n159 86.7903
R548 VSS.n2188 VSS.n2187 86.7903
R549 VSS.n2182 VSS.n166 86.7903
R550 VSS.t5 VSS.n197 85.0843
R551 VSS.n1028 VSS.n1027 82.5693
R552 VSS.n2295 VSS.n2294 80.858
R553 VSS.n778 VSS.n774 80.0913
R554 VSS.n838 VSS.n318 80.0913
R555 VSS.n1630 VSS.n1629 80.0913
R556 VSS.n1713 VSS.n259 80.0913
R557 VSS.t1 VSS.t23 78.4806
R558 VSS.n1886 VSS.n1885 76.183
R559 VSS.n992 VSS.n703 75.6886
R560 VSS.n1207 VSS.n577 75.3628
R561 VSS.n1335 VSS.n523 75.3628
R562 VSS.n1496 VSS.n470 75.3628
R563 VSS.n1430 VSS.n327 75.3628
R564 VSS.n2343 VSS.n17 75.3628
R565 VSS.n1091 VSS.n1090 71.4377
R566 VSS.n228 VSS.n223 70.8914
R567 VSS.n2294 VSS.n44 69.8676
R568 VSS.n2128 VSS.n2127 67.4011
R569 VSS.n1090 VSS.n620 64.3725
R570 VSS.n1149 VSS.n1148 62.8024
R571 VSS.n1277 VSS.n1276 62.8024
R572 VSS.n1405 VSS.n1404 62.8024
R573 VSS.n1425 VSS.n425 62.8024
R574 VSS.n1572 VSS.n346 62.8024
R575 VSS.n1906 VSS.n1905 57.4122
R576 VSS.n2012 VSS.n63 51.9206
R577 VSS.n2209 VSS.t19 51.2434
R578 VSS.n1133 VSS.t2 49.457
R579 VSS.n1261 VSS.t15 49.457
R580 VSS.n1389 VSS.t7 49.457
R581 VSS.n1447 VSS.t9 49.457
R582 VSS.n1589 VSS.t13 49.457
R583 VSS.t0 VSS.n44 49.457
R584 VSS.n2236 VSS.n63 47.9268
R585 VSS.n2103 VSS.n2102 46.1653
R586 VSS.n2181 VSS.n169 44.3187
R587 VSS.n2078 VSS.n2077 43.857
R588 VSS.n1907 VSS.t11 43.4337
R589 VSS.n2078 VSS.n165 42.9337
R590 VSS.n2293 VSS.n46 36.7314
R591 VSS.n1091 VSS.n619 35.3266
R592 VSS.n2029 VSS.n207 34.7841
R593 VSS.n1952 VSS.n1951 31.4521
R594 VSS.n709 VSS.n197 24.4653
R595 VSS.n1948 VSS.n228 22.9652
R596 VSS.n2208 VSS.t3 21.6979
R597 VSS.n142 VSS.n136 20.9682
R598 VSS.n2061 VSS.n198 20.7673
R599 VSS.t22 VSS.t19 20.313
R600 VSS.n2128 VSS.n151 19.3897
R601 VSS.n1093 VSS.n617 19.3426
R602 VSS.n1952 VSS.t11 18.9713
R603 VSS.n2103 VSS.t3 18.9281
R604 VSS.n2088 VSS.n179 18.4216
R605 VSS.n2093 VSS.n2092 18.4216
R606 VSS.n2097 VSS.n2096 18.4216
R607 VSS.n2099 VSS.n175 18.4216
R608 VSS.n2107 VSS.n175 18.4216
R609 VSS.n2111 VSS.n2109 18.4216
R610 VSS.n2115 VSS.n173 18.4216
R611 VSS.n2118 VSS.n2117 18.4216
R612 VSS.n2030 VSS.n1984 18.4216
R613 VSS.n2026 VSS.n1984 18.4216
R614 VSS.n2026 VSS.n1987 18.4216
R615 VSS.n2022 VSS.n1987 18.4216
R616 VSS.n2022 VSS.n1990 18.4216
R617 VSS.n2018 VSS.n1990 18.4216
R618 VSS.n2018 VSS.n1992 18.4216
R619 VSS.n2014 VSS.n1992 18.4216
R620 VSS.n2014 VSS.n2011 18.4216
R621 VSS.n2009 VSS.n1994 18.4216
R622 VSS.n2005 VSS.n2004 18.4216
R623 VSS.n2002 VSS.n1999 18.4216
R624 VSS.n1727 VSS.n284 18.4216
R625 VSS.n1723 VSS.n284 18.4216
R626 VSS.n1723 VSS.n1687 18.4216
R627 VSS.n1719 VSS.n1687 18.4216
R628 VSS.n1719 VSS.n1689 18.4216
R629 VSS.n1715 VSS.n1689 18.4216
R630 VSS.n1715 VSS.n1712 18.4216
R631 VSS.n1712 VSS.n1711 18.4216
R632 VSS.n1711 VSS.n1691 18.4216
R633 VSS.n1707 VSS.n1691 18.4216
R634 VSS.n1707 VSS.n1694 18.4216
R635 VSS.n1703 VSS.n1694 18.4216
R636 VSS.n1703 VSS.n1701 18.4216
R637 VSS.n1698 VSS.n1697 18.4216
R638 VSS.n1644 VSS.n308 18.4216
R639 VSS.n1640 VSS.n308 18.4216
R640 VSS.n1640 VSS.n313 18.4216
R641 VSS.n1636 VSS.n313 18.4216
R642 VSS.n1636 VSS.n315 18.4216
R643 VSS.n1632 VSS.n315 18.4216
R644 VSS.n1632 VSS.n317 18.4216
R645 VSS.n1627 VSS.n317 18.4216
R646 VSS.n1627 VSS.n320 18.4216
R647 VSS.n1623 VSS.n320 18.4216
R648 VSS.n1623 VSS.n322 18.4216
R649 VSS.n1619 VSS.n322 18.4216
R650 VSS.n1619 VSS.n324 18.4216
R651 VSS.n1615 VSS.n1614 18.4216
R652 VSS.n875 VSS.n833 18.4216
R653 VSS.n871 VSS.n833 18.4216
R654 VSS.n871 VSS.n835 18.4216
R655 VSS.n867 VSS.n835 18.4216
R656 VSS.n867 VSS.n837 18.4216
R657 VSS.n863 VSS.n837 18.4216
R658 VSS.n863 VSS.n839 18.4216
R659 VSS.n859 VSS.n839 18.4216
R660 VSS.n859 VSS.n841 18.4216
R661 VSS.n855 VSS.n841 18.4216
R662 VSS.n855 VSS.n843 18.4216
R663 VSS.n851 VSS.n843 18.4216
R664 VSS.n851 VSS.n849 18.4216
R665 VSS.n846 VSS.n845 18.4216
R666 VSS.n812 VSS.n769 18.4216
R667 VSS.n808 VSS.n769 18.4216
R668 VSS.n808 VSS.n771 18.4216
R669 VSS.n804 VSS.n771 18.4216
R670 VSS.n804 VSS.n773 18.4216
R671 VSS.n800 VSS.n773 18.4216
R672 VSS.n800 VSS.n775 18.4216
R673 VSS.n796 VSS.n775 18.4216
R674 VSS.n796 VSS.n777 18.4216
R675 VSS.n792 VSS.n777 18.4216
R676 VSS.n792 VSS.n780 18.4216
R677 VSS.n788 VSS.n780 18.4216
R678 VSS.n788 VSS.n786 18.4216
R679 VSS.n783 VSS.n782 18.4216
R680 VSS.n1026 VSS.n995 18.4216
R681 VSS.n1022 VSS.n1021 18.4216
R682 VSS.n1018 VSS.n1017 18.4216
R683 VSS.n1014 VSS.n1013 18.4216
R684 VSS.n1010 VSS.n1009 18.4216
R685 VSS.n1006 VSS.n1005 18.4216
R686 VSS.n1002 VSS.n1001 18.4216
R687 VSS.n998 VSS.n997 18.4216
R688 VSS.n671 VSS.n670 18.4216
R689 VSS.n667 VSS.n666 18.4216
R690 VSS.n664 VSS.n626 18.4216
R691 VSS.n660 VSS.n658 18.4216
R692 VSS.n656 VSS.n628 18.4216
R693 VSS.n652 VSS.n650 18.4216
R694 VSS.n648 VSS.n630 18.4216
R695 VSS.n644 VSS.n642 18.4216
R696 VSS.n642 VSS.n641 18.4216
R697 VSS.n638 VSS.n637 18.4216
R698 VSS.n635 VSS.n617 18.4216
R699 VSS.n1206 VSS.n589 18.4216
R700 VSS.n1202 VSS.n1201 18.4216
R701 VSS.n1198 VSS.n1197 18.4216
R702 VSS.n1194 VSS.n1193 18.4216
R703 VSS.n1190 VSS.n1189 18.4216
R704 VSS.n1186 VSS.n1185 18.4216
R705 VSS.n1182 VSS.n1181 18.4216
R706 VSS.n1209 VSS.n576 18.4216
R707 VSS.n1218 VSS.n573 18.4216
R708 VSS.n1218 VSS.n574 18.4216
R709 VSS.n1214 VSS.n1213 18.4216
R710 VSS.n1334 VSS.n535 18.4216
R711 VSS.n1330 VSS.n1329 18.4216
R712 VSS.n1326 VSS.n1325 18.4216
R713 VSS.n1322 VSS.n1321 18.4216
R714 VSS.n1318 VSS.n1317 18.4216
R715 VSS.n1314 VSS.n1313 18.4216
R716 VSS.n1310 VSS.n1309 18.4216
R717 VSS.n1337 VSS.n522 18.4216
R718 VSS.n1346 VSS.n519 18.4216
R719 VSS.n1346 VSS.n520 18.4216
R720 VSS.n1342 VSS.n1341 18.4216
R721 VSS.n1495 VSS.n482 18.4216
R722 VSS.n1491 VSS.n1490 18.4216
R723 VSS.n1487 VSS.n1486 18.4216
R724 VSS.n1483 VSS.n1482 18.4216
R725 VSS.n1479 VSS.n1478 18.4216
R726 VSS.n1475 VSS.n1474 18.4216
R727 VSS.n1471 VSS.n1470 18.4216
R728 VSS.n1498 VSS.n469 18.4216
R729 VSS.n1507 VSS.n466 18.4216
R730 VSS.n1507 VSS.n467 18.4216
R731 VSS.n1503 VSS.n1502 18.4216
R732 VSS.n383 VSS.n381 18.4216
R733 VSS.n387 VSS.n380 18.4216
R734 VSS.n391 VSS.n389 18.4216
R735 VSS.n395 VSS.n378 18.4216
R736 VSS.n399 VSS.n397 18.4216
R737 VSS.n403 VSS.n376 18.4216
R738 VSS.n407 VSS.n405 18.4216
R739 VSS.n411 VSS.n374 18.4216
R740 VSS.n414 VSS.n413 18.4216
R741 VSS.n415 VSS.n414 18.4216
R742 VSS.n419 VSS.n418 18.4216
R743 VSS.n2342 VSS.n29 18.4216
R744 VSS.n2338 VSS.n2337 18.4216
R745 VSS.n2334 VSS.n2333 18.4216
R746 VSS.n2330 VSS.n2329 18.4216
R747 VSS.n2326 VSS.n2325 18.4216
R748 VSS.n2322 VSS.n2321 18.4216
R749 VSS.n2318 VSS.n2317 18.4216
R750 VSS.n2345 VSS.n16 18.4216
R751 VSS.n2354 VSS.n13 18.4216
R752 VSS.n2354 VSS.n14 18.4216
R753 VSS.n2350 VSS.n2349 18.4216
R754 VSS.n737 VSS.n723 18.4216
R755 VSS.n737 VSS.n725 18.4216
R756 VSS.n733 VSS.n725 18.4216
R757 VSS.n733 VSS.n727 18.4216
R758 VSS.n729 VSS.n727 18.4216
R759 VSS.n729 VSS.n683 18.4216
R760 VSS.n1047 VSS.n683 18.4216
R761 VSS.n1047 VSS.n681 18.4216
R762 VSS.n1051 VSS.n681 18.4216
R763 VSS.n1051 VSS.n679 18.4216
R764 VSS.n1056 VSS.n679 18.4216
R765 VSS.n1056 VSS.n677 18.4216
R766 VSS.n1060 VSS.n677 18.4216
R767 VSS.n1063 VSS.n1062 18.4216
R768 VSS.n762 VSS.n761 18.4216
R769 VSS.n759 VSS.n742 18.4216
R770 VSS.n755 VSS.n754 18.4216
R771 VSS.n752 VSS.n745 18.4216
R772 VSS.n748 VSS.n745 18.4216
R773 VSS.n748 VSS.n687 18.4216
R774 VSS.n1042 VSS.n687 18.4216
R775 VSS.n1042 VSS.n688 18.4216
R776 VSS.n1038 VSS.n688 18.4216
R777 VSS.n1038 VSS.n691 18.4216
R778 VSS.n1034 VSS.n691 18.4216
R779 VSS.n1034 VSS.n693 18.4216
R780 VSS.n1030 VSS.n693 18.4216
R781 VSS.n1030 VSS.n695 18.4216
R782 VSS.n993 VSS.n702 18.4216
R783 VSS.n989 VSS.n702 18.4216
R784 VSS.n989 VSS.n705 18.4216
R785 VSS.n985 VSS.n705 18.4216
R786 VSS.n985 VSS.n708 18.4216
R787 VSS.n981 VSS.n708 18.4216
R788 VSS.n981 VSS.n710 18.4216
R789 VSS.n977 VSS.n710 18.4216
R790 VSS.n977 VSS.n712 18.4216
R791 VSS.n974 VSS.n713 18.4216
R792 VSS.n970 VSS.n969 18.4216
R793 VSS.n967 VSS.n717 18.4216
R794 VSS.n963 VSS.n962 18.4216
R795 VSS.n954 VSS.n815 18.4216
R796 VSS.n950 VSS.n949 18.4216
R797 VSS.n947 VSS.n818 18.4216
R798 VSS.n943 VSS.n942 18.4216
R799 VSS.n942 VSS.n821 18.4216
R800 VSS.n939 VSS.n822 18.4216
R801 VSS.n935 VSS.n934 18.4216
R802 VSS.n932 VSS.n827 18.4216
R803 VSS.n928 VSS.n927 18.4216
R804 VSS.n919 VSS.n878 18.4216
R805 VSS.n915 VSS.n914 18.4216
R806 VSS.n912 VSS.n881 18.4216
R807 VSS.n908 VSS.n907 18.4216
R808 VSS.n907 VSS.n884 18.4216
R809 VSS.n904 VSS.n885 18.4216
R810 VSS.n900 VSS.n899 18.4216
R811 VSS.n896 VSS.n895 18.4216
R812 VSS.n892 VSS.n891 18.4216
R813 VSS.n300 VSS.n299 18.4216
R814 VSS.n304 VSS.n297 18.4216
R815 VSS.n1648 VSS.n290 18.4216
R816 VSS.n1653 VSS.n288 18.4216
R817 VSS.n1653 VSS.n287 18.4216
R818 VSS.n1657 VSS.n1656 18.4216
R819 VSS.n1661 VSS.n1660 18.4216
R820 VSS.n1665 VSS.n1664 18.4216
R821 VSS.n1669 VSS.n1668 18.4216
R822 VSS.n1680 VSS.n1679 18.4216
R823 VSS.n1676 VSS.n1675 18.4216
R824 VSS.n1731 VSS.n274 18.4216
R825 VSS.n1736 VSS.n272 18.4216
R826 VSS.n1736 VSS.n271 18.4216
R827 VSS.n1741 VSS.n1739 18.4216
R828 VSS.n1745 VSS.n269 18.4216
R829 VSS.n1749 VSS.n1747 18.4216
R830 VSS.n1753 VSS.n267 18.4216
R831 VSS.n1978 VSS.n1977 18.4216
R832 VSS.n1975 VSS.n220 18.4216
R833 VSS.n1971 VSS.n1970 18.4216
R834 VSS.n1968 VSS.n1954 18.4216
R835 VSS.n1964 VSS.n1963 18.4216
R836 VSS.n1961 VSS.n1958 18.4216
R837 VSS.n2059 VSS.n213 18.4216
R838 VSS.n2059 VSS.n214 18.4216
R839 VSS.n2055 VSS.n2054 18.4216
R840 VSS.n2044 VSS.n2043 18.4216
R841 VSS.n2040 VSS.n2039 18.4216
R842 VSS.n2036 VSS.n2035 18.4216
R843 VSS.n2035 VSS.n2034 18.4216
R844 VSS.n2063 VSS.n195 18.4216
R845 VSS.n2063 VSS.n193 18.4216
R846 VSS.n2067 VSS.n193 18.4216
R847 VSS.n2067 VSS.n191 18.4216
R848 VSS.n2071 VSS.n191 18.4216
R849 VSS.n2071 VSS.n189 18.4216
R850 VSS.n2075 VSS.n189 18.4216
R851 VSS.n2075 VSS.n187 18.4216
R852 VSS.n2082 VSS.n187 18.4216
R853 VSS.n2082 VSS.n185 18.4216
R854 VSS.n1759 VSS.n265 18.4216
R855 VSS.n1763 VSS.n265 18.4216
R856 VSS.n1763 VSS.n263 18.4216
R857 VSS.n1767 VSS.n263 18.4216
R858 VSS.n1767 VSS.n261 18.4216
R859 VSS.n1771 VSS.n261 18.4216
R860 VSS.n1771 VSS.n258 18.4216
R861 VSS.n1776 VSS.n258 18.4216
R862 VSS.n1776 VSS.n256 18.4216
R863 VSS.n1780 VSS.n256 18.4216
R864 VSS.n1780 VSS.n254 18.4216
R865 VSS.n1784 VSS.n254 18.4216
R866 VSS.n1784 VSS.n252 18.4216
R867 VSS.n1788 VSS.n252 18.4216
R868 VSS.n1788 VSS.n250 18.4216
R869 VSS.n1792 VSS.n250 18.4216
R870 VSS.n1836 VSS.n246 18.4216
R871 VSS.n1840 VSS.n246 18.4216
R872 VSS.n1840 VSS.n244 18.4216
R873 VSS.n1844 VSS.n244 18.4216
R874 VSS.n1844 VSS.n241 18.4216
R875 VSS.n1849 VSS.n241 18.4216
R876 VSS.n1849 VSS.n238 18.4216
R877 VSS.n1884 VSS.n238 18.4216
R878 VSS.n1884 VSS.n239 18.4216
R879 VSS.n1880 VSS.n239 18.4216
R880 VSS.n1880 VSS.n1853 18.4216
R881 VSS.n1876 VSS.n1853 18.4216
R882 VSS.n1876 VSS.n1855 18.4216
R883 VSS.n1872 VSS.n1855 18.4216
R884 VSS.n1872 VSS.n1857 18.4216
R885 VSS.n1868 VSS.n1857 18.4216
R886 VSS.n1868 VSS.n1859 18.4216
R887 VSS.n1864 VSS.n1859 18.4216
R888 VSS.n1864 VSS.n1861 18.4216
R889 VSS.n1861 VSS.n48 18.4216
R890 VSS.n2291 VSS.n48 18.4216
R891 VSS.n1089 VSS.n622 18.4216
R892 VSS.n1085 VSS.n622 18.4216
R893 VSS.n1085 VSS.n1069 18.4216
R894 VSS.n1081 VSS.n1069 18.4216
R895 VSS.n1081 VSS.n1072 18.4216
R896 VSS.n1077 VSS.n1072 18.4216
R897 VSS.n1077 VSS.n1074 18.4216
R898 VSS.n1074 VSS.n603 18.4216
R899 VSS.n1134 VSS.n603 18.4216
R900 VSS.n1134 VSS.n601 18.4216
R901 VSS.n1138 VSS.n601 18.4216
R902 VSS.n1138 VSS.n599 18.4216
R903 VSS.n1142 VSS.n599 18.4216
R904 VSS.n1142 VSS.n597 18.4216
R905 VSS.n1147 VSS.n597 18.4216
R906 VSS.n1147 VSS.n593 18.4216
R907 VSS.n1152 VSS.n593 18.4216
R908 VSS.n1153 VSS.n1152 18.4216
R909 VSS.n1177 VSS.n1156 18.4216
R910 VSS.n1173 VSS.n1156 18.4216
R911 VSS.n1173 VSS.n1158 18.4216
R912 VSS.n1169 VSS.n1158 18.4216
R913 VSS.n1169 VSS.n1160 18.4216
R914 VSS.n1165 VSS.n1160 18.4216
R915 VSS.n1165 VSS.n1162 18.4216
R916 VSS.n1162 VSS.n549 18.4216
R917 VSS.n1262 VSS.n549 18.4216
R918 VSS.n1262 VSS.n547 18.4216
R919 VSS.n1266 VSS.n547 18.4216
R920 VSS.n1266 VSS.n545 18.4216
R921 VSS.n1270 VSS.n545 18.4216
R922 VSS.n1270 VSS.n543 18.4216
R923 VSS.n1275 VSS.n543 18.4216
R924 VSS.n1275 VSS.n539 18.4216
R925 VSS.n1280 VSS.n539 18.4216
R926 VSS.n1281 VSS.n1280 18.4216
R927 VSS.n1305 VSS.n1284 18.4216
R928 VSS.n1301 VSS.n1284 18.4216
R929 VSS.n1301 VSS.n1286 18.4216
R930 VSS.n1297 VSS.n1286 18.4216
R931 VSS.n1297 VSS.n1288 18.4216
R932 VSS.n1293 VSS.n1288 18.4216
R933 VSS.n1293 VSS.n1290 18.4216
R934 VSS.n1290 VSS.n496 18.4216
R935 VSS.n1390 VSS.n496 18.4216
R936 VSS.n1390 VSS.n494 18.4216
R937 VSS.n1394 VSS.n494 18.4216
R938 VSS.n1394 VSS.n492 18.4216
R939 VSS.n1398 VSS.n492 18.4216
R940 VSS.n1398 VSS.n490 18.4216
R941 VSS.n1403 VSS.n490 18.4216
R942 VSS.n1403 VSS.n486 18.4216
R943 VSS.n1408 VSS.n486 18.4216
R944 VSS.n1409 VSS.n1408 18.4216
R945 VSS.n1466 VSS.n1412 18.4216
R946 VSS.n1462 VSS.n1412 18.4216
R947 VSS.n1462 VSS.n1414 18.4216
R948 VSS.n1458 VSS.n1414 18.4216
R949 VSS.n1458 VSS.n1416 18.4216
R950 VSS.n1454 VSS.n1416 18.4216
R951 VSS.n1454 VSS.n1418 18.4216
R952 VSS.n1450 VSS.n1418 18.4216
R953 VSS.n1450 VSS.n1420 18.4216
R954 VSS.n1445 VSS.n1420 18.4216
R955 VSS.n1445 VSS.n1422 18.4216
R956 VSS.n1441 VSS.n1422 18.4216
R957 VSS.n1441 VSS.n1424 18.4216
R958 VSS.n1437 VSS.n1424 18.4216
R959 VSS.n1437 VSS.n1426 18.4216
R960 VSS.n1433 VSS.n1426 18.4216
R961 VSS.n1433 VSS.n1428 18.4216
R962 VSS.n1429 VSS.n1428 18.4216
R963 VSS.n1608 VSS.n332 18.4216
R964 VSS.n1604 VSS.n332 18.4216
R965 VSS.n1604 VSS.n334 18.4216
R966 VSS.n1600 VSS.n334 18.4216
R967 VSS.n1600 VSS.n336 18.4216
R968 VSS.n1596 VSS.n336 18.4216
R969 VSS.n1596 VSS.n338 18.4216
R970 VSS.n1592 VSS.n338 18.4216
R971 VSS.n1592 VSS.n340 18.4216
R972 VSS.n1587 VSS.n340 18.4216
R973 VSS.n1587 VSS.n343 18.4216
R974 VSS.n1583 VSS.n343 18.4216
R975 VSS.n1583 VSS.n345 18.4216
R976 VSS.n1579 VSS.n345 18.4216
R977 VSS.n1579 VSS.n347 18.4216
R978 VSS.n1575 VSS.n347 18.4216
R979 VSS.n1575 VSS.n350 18.4216
R980 VSS.n350 VSS.n349 18.4216
R981 VSS.n2313 VSS.n34 18.4216
R982 VSS.n2309 VSS.n34 18.4216
R983 VSS.n2309 VSS.n36 18.4216
R984 VSS.n2305 VSS.n36 18.4216
R985 VSS.n2305 VSS.n38 18.4216
R986 VSS.n2301 VSS.n38 18.4216
R987 VSS.n2301 VSS.n40 18.4216
R988 VSS.n2297 VSS.n40 18.4216
R989 VSS.n2297 VSS.n42 18.4216
R990 VSS.n1799 VSS.n42 18.4216
R991 VSS.n1801 VSS.n1799 18.4216
R992 VSS.n1805 VSS.n1797 18.4216
R993 VSS.n1808 VSS.n1807 18.4216
R994 VSS.n1812 VSS.n1811 18.4216
R995 VSS.n1830 VSS.n1829 18.4216
R996 VSS.n1827 VSS.n1818 18.4216
R997 VSS.n1823 VSS.n1822 18.4216
R998 VSS.n1908 VSS.n233 18.4216
R999 VSS.n1908 VSS.n230 18.4216
R1000 VSS.n1946 VSS.n230 18.4216
R1001 VSS.n1946 VSS.n231 18.4216
R1002 VSS.n1942 VSS.n231 18.4216
R1003 VSS.n1942 VSS.n1912 18.4216
R1004 VSS.n1925 VSS.n1912 18.4216
R1005 VSS.n1932 VSS.n1925 18.4216
R1006 VSS.n1932 VSS.n1928 18.4216
R1007 VSS.n1928 VSS.n64 18.4216
R1008 VSS.n2235 VSS.n64 18.4216
R1009 VSS.n2231 VSS.n125 18.4216
R1010 VSS.n2224 VSS.n125 18.4216
R1011 VSS.n2224 VSS.n131 18.4216
R1012 VSS.n2220 VSS.n131 18.4216
R1013 VSS.n2220 VSS.n133 18.4216
R1014 VSS.n204 VSS.n133 18.4216
R1015 VSS.n204 VSS.n201 18.4216
R1016 VSS.n2207 VSS.n145 18.4216
R1017 VSS.n2207 VSS.n146 18.4216
R1018 VSS.n2203 VSS.n146 18.4216
R1019 VSS.n2203 VSS.n149 18.4216
R1020 VSS.n160 VSS.n149 18.4216
R1021 VSS.n2193 VSS.n160 18.4216
R1022 VSS.n2193 VSS.n161 18.4216
R1023 VSS.n2189 VSS.n161 18.4216
R1024 VSS.n2189 VSS.n164 18.4216
R1025 VSS.n2180 VSS.n164 18.4216
R1026 VSS.n2174 VSS.n2173 18.4216
R1027 VSS.n2170 VSS.n2169 18.4216
R1028 VSS.n2167 VSS.n2125 18.4216
R1029 VSS.n2163 VSS.n2161 18.4216
R1030 VSS.n2159 VSS.n2129 18.4216
R1031 VSS.n2155 VSS.n2153 18.4216
R1032 VSS.n2151 VSS.n2131 18.4216
R1033 VSS.n2147 VSS.n2145 18.4216
R1034 VSS.n2143 VSS.n2133 18.4216
R1035 VSS.n2139 VSS.n2137 18.4216
R1036 VSS.n1093 VSS.n615 18.4216
R1037 VSS.n1097 VSS.n615 18.4216
R1038 VSS.n1097 VSS.n613 18.4216
R1039 VSS.n1101 VSS.n613 18.4216
R1040 VSS.n1101 VSS.n611 18.4216
R1041 VSS.n1105 VSS.n611 18.4216
R1042 VSS.n1105 VSS.n608 18.4216
R1043 VSS.n1129 VSS.n608 18.4216
R1044 VSS.n1129 VSS.n609 18.4216
R1045 VSS.n1125 VSS.n609 18.4216
R1046 VSS.n1125 VSS.n1109 18.4216
R1047 VSS.n1121 VSS.n1109 18.4216
R1048 VSS.n1121 VSS.n1111 18.4216
R1049 VSS.n1117 VSS.n1111 18.4216
R1050 VSS.n1117 VSS.n1112 18.4216
R1051 VSS.n1113 VSS.n1112 18.4216
R1052 VSS.n1113 VSS.n566 18.4216
R1053 VSS.n1221 VSS.n566 18.4216
R1054 VSS.n564 VSS.n561 18.4216
R1055 VSS.n1225 VSS.n561 18.4216
R1056 VSS.n1225 VSS.n559 18.4216
R1057 VSS.n1229 VSS.n559 18.4216
R1058 VSS.n1229 VSS.n557 18.4216
R1059 VSS.n1233 VSS.n557 18.4216
R1060 VSS.n1233 VSS.n554 18.4216
R1061 VSS.n1257 VSS.n554 18.4216
R1062 VSS.n1257 VSS.n555 18.4216
R1063 VSS.n1253 VSS.n555 18.4216
R1064 VSS.n1253 VSS.n1237 18.4216
R1065 VSS.n1249 VSS.n1237 18.4216
R1066 VSS.n1249 VSS.n1239 18.4216
R1067 VSS.n1245 VSS.n1239 18.4216
R1068 VSS.n1245 VSS.n1240 18.4216
R1069 VSS.n1241 VSS.n1240 18.4216
R1070 VSS.n1241 VSS.n512 18.4216
R1071 VSS.n1349 VSS.n512 18.4216
R1072 VSS.n510 VSS.n507 18.4216
R1073 VSS.n1353 VSS.n507 18.4216
R1074 VSS.n1353 VSS.n505 18.4216
R1075 VSS.n1357 VSS.n505 18.4216
R1076 VSS.n1357 VSS.n503 18.4216
R1077 VSS.n1361 VSS.n503 18.4216
R1078 VSS.n1361 VSS.n500 18.4216
R1079 VSS.n1385 VSS.n500 18.4216
R1080 VSS.n1385 VSS.n501 18.4216
R1081 VSS.n1381 VSS.n501 18.4216
R1082 VSS.n1381 VSS.n1365 18.4216
R1083 VSS.n1377 VSS.n1365 18.4216
R1084 VSS.n1377 VSS.n1367 18.4216
R1085 VSS.n1373 VSS.n1367 18.4216
R1086 VSS.n1373 VSS.n1368 18.4216
R1087 VSS.n1369 VSS.n1368 18.4216
R1088 VSS.n1369 VSS.n442 18.4216
R1089 VSS.n1510 VSS.n442 18.4216
R1090 VSS.n460 VSS.n441 18.4216
R1091 VSS.n460 VSS.n459 18.4216
R1092 VSS.n459 VSS.n446 18.4216
R1093 VSS.n455 VSS.n446 18.4216
R1094 VSS.n455 VSS.n448 18.4216
R1095 VSS.n451 VSS.n448 18.4216
R1096 VSS.n451 VSS.n434 18.4216
R1097 VSS.n1515 VSS.n434 18.4216
R1098 VSS.n1515 VSS.n432 18.4216
R1099 VSS.n1519 VSS.n432 18.4216
R1100 VSS.n1519 VSS.n430 18.4216
R1101 VSS.n1523 VSS.n430 18.4216
R1102 VSS.n1523 VSS.n428 18.4216
R1103 VSS.n1528 VSS.n428 18.4216
R1104 VSS.n1528 VSS.n426 18.4216
R1105 VSS.n1532 VSS.n426 18.4216
R1106 VSS.n1532 VSS.n424 18.4216
R1107 VSS.n1536 VSS.n424 18.4216
R1108 VSS.n1538 VSS.n366 18.4216
R1109 VSS.n1542 VSS.n366 18.4216
R1110 VSS.n1542 VSS.n364 18.4216
R1111 VSS.n1546 VSS.n364 18.4216
R1112 VSS.n1546 VSS.n362 18.4216
R1113 VSS.n1550 VSS.n362 18.4216
R1114 VSS.n1550 VSS.n360 18.4216
R1115 VSS.n1554 VSS.n360 18.4216
R1116 VSS.n1554 VSS.n358 18.4216
R1117 VSS.n1558 VSS.n358 18.4216
R1118 VSS.n1558 VSS.n356 18.4216
R1119 VSS.n1562 VSS.n356 18.4216
R1120 VSS.n1562 VSS.n354 18.4216
R1121 VSS.n1566 VSS.n354 18.4216
R1122 VSS.n1566 VSS.n352 18.4216
R1123 VSS.n1570 VSS.n352 18.4216
R1124 VSS.n1570 VSS.n6 18.4216
R1125 VSS.n2357 VSS.n6 18.4216
R1126 VSS.n2253 VSS.n5 18.4216
R1127 VSS.n2256 VSS.n2253 18.4216
R1128 VSS.n2256 VSS.n2252 18.4216
R1129 VSS.n2260 VSS.n2252 18.4216
R1130 VSS.n2260 VSS.n2250 18.4216
R1131 VSS.n2264 VSS.n2250 18.4216
R1132 VSS.n2264 VSS.n2248 18.4216
R1133 VSS.n2269 VSS.n2247 18.4216
R1134 VSS.n2275 VSS.n2273 18.4216
R1135 VSS.n2279 VSS.n2245 18.4216
R1136 VSS.n2282 VSS.n2281 18.4216
R1137 VSS.n2286 VSS.n2285 18.4216
R1138 VSS.n1892 VSS.n1890 18.4216
R1139 VSS.n1895 VSS.n1894 18.4216
R1140 VSS.n1897 VSS.n1887 18.4216
R1141 VSS.n1902 VSS.n224 18.4216
R1142 VSS.n1950 VSS.n224 18.4216
R1143 VSS.n1950 VSS.n1949 18.4216
R1144 VSS.n1949 VSS.n225 18.4216
R1145 VSS.n1916 VSS.n225 18.4216
R1146 VSS.n1939 VSS.n1916 18.4216
R1147 VSS.n1939 VSS.n1917 18.4216
R1148 VSS.n1935 VSS.n1917 18.4216
R1149 VSS.n1935 VSS.n1921 18.4216
R1150 VSS.n1921 VSS.n60 18.4216
R1151 VSS.n2238 VSS.n60 18.4216
R1152 VSS.n2228 VSS.n59 18.4216
R1153 VSS.n2228 VSS.n2227 18.4216
R1154 VSS.n2227 VSS.n128 18.4216
R1155 VSS.n137 VSS.n128 18.4216
R1156 VSS.n2217 VSS.n137 18.4216
R1157 VSS.n2217 VSS.n138 18.4216
R1158 VSS.n2213 VSS.n138 18.4216
R1159 VSS.n2211 VSS.n2210 18.4216
R1160 VSS.n2210 VSS.n143 18.4216
R1161 VSS.n152 VSS.n143 18.4216
R1162 VSS.n2200 VSS.n152 18.4216
R1163 VSS.n2200 VSS.n153 18.4216
R1164 VSS.n2196 VSS.n153 18.4216
R1165 VSS.n2196 VSS.n157 18.4216
R1166 VSS.n167 VSS.n157 18.4216
R1167 VSS.n2186 VSS.n167 18.4216
R1168 VSS.n2186 VSS.n2183 18.4216
R1169 VSS.n121 VSS.n120 18.4216
R1170 VSS.n118 VSS.n68 18.4216
R1171 VSS.n114 VSS.n112 18.4216
R1172 VSS.n110 VSS.n70 18.4216
R1173 VSS.n106 VSS.n104 18.4216
R1174 VSS.n102 VSS.n72 18.4216
R1175 VSS.n98 VSS.n96 18.4216
R1176 VSS.n94 VSS.n74 18.4216
R1177 VSS.n90 VSS.n88 18.4216
R1178 VSS.n86 VSS.n79 18.4216
R1179 VSS.n82 VSS.n80 18.4216
R1180 VSS.n764 VSS.n723 17.8689
R1181 VSS.n2183 VSS.n168 17.8689
R1182 VSS.n185 VSS.n181 16.3952
R1183 VSS.n1044 VSS.n1043 15.291
R1184 VSS.n2104 VSS.n2103 12.5416
R1185 VSS.n1089 VSS.n621 12.5268
R1186 VSS.n1177 VSS.n588 12.5268
R1187 VSS.n1305 VSS.n534 12.5268
R1188 VSS.n1466 VSS.n481 12.5268
R1189 VSS.n1608 VSS.n328 12.5268
R1190 VSS.n2313 VSS.n28 12.5268
R1191 VSS.n1832 VSS.n248 12.5268
R1192 VSS.n2231 VSS.n65 12.5268
R1193 VSS.n1131 VSS.t17 12.3005
R1194 VSS.n1259 VSS.t16 12.3005
R1195 VSS.n1387 VSS.t8 12.3005
R1196 VSS.n436 VSS.t10 12.3005
R1197 VSS.n341 VSS.t14 12.3005
R1198 VSS.n227 VSS.t12 12.3005
R1199 VSS.n43 VSS.t18 12.3005
R1200 VSS.n994 VSS.n993 11.4216
R1201 VSS.n956 VSS.n720 11.4216
R1202 VSS.n921 VSS.n830 11.4216
R1203 VSS.n309 VSS.n307 11.4216
R1204 VSS.n1683 VSS.n283 11.4216
R1205 VSS.n1980 VSS.n217 11.4216
R1206 VSS.n2049 VSS.n2048 11.4216
R1207 VSS.n567 VSS.n564 11.4216
R1208 VSS.n513 VSS.n510 11.4216
R1209 VSS.n443 VSS.n441 11.4216
R1210 VSS.n1538 VSS.n368 11.4216
R1211 VSS.n7 VSS.n5 11.4216
R1212 VSS.n53 VSS.n49 11.4216
R1213 VSS.n61 VSS.n59 11.4216
R1214 VSS.n182 VSS.t6 11.2214
R1215 VSS.n1207 VSS.n587 10.9908
R1216 VSS.n1335 VSS.n533 10.9908
R1217 VSS.n1496 VSS.n480 10.9908
R1218 VSS.n327 VSS.n323 10.9908
R1219 VSS.n2343 VSS.n27 10.9908
R1220 VSS.n1027 VSS.n587 10.7039
R1221 VSS.n228 VSS.n227 10.4005
R1222 VSS.n183 VSS.n180 10.4005
R1223 VSS.n182 VSS.n180 10.4005
R1224 VSS.n1903 VSS.n1887 10.3636
R1225 VSS.n1822 VSS.n1821 10.3596
R1226 VSS.n2012 VSS.n126 9.98514
R1227 VSS.n994 VSS.n695 9.94787
R1228 VSS.n960 VSS.n720 9.94787
R1229 VSS.n925 VSS.n830 9.94787
R1230 VSS.n887 VSS.n307 9.94787
R1231 VSS.n1672 VSS.n283 9.94787
R1232 VSS.n1755 VSS.n217 9.94787
R1233 VSS.n2050 VSS.n2049 9.94787
R1234 VSS.n1221 VSS.n567 9.94787
R1235 VSS.n1349 VSS.n513 9.94787
R1236 VSS.n1510 VSS.n443 9.94787
R1237 VSS.n1536 VSS.n368 9.94787
R1238 VSS.n2357 VSS.n7 9.94787
R1239 VSS.n2288 VSS.n49 9.94787
R1240 VSS.n2238 VSS.n61 9.94787
R1241 VSS.n1153 VSS.n588 8.84261
R1242 VSS.n1281 VSS.n534 8.84261
R1243 VSS.n1409 VSS.n481 8.84261
R1244 VSS.n1429 VSS.n328 8.84261
R1245 VSS.n349 VSS.n28 8.84261
R1246 VSS.n1814 VSS.n248 8.84261
R1247 VSS.n2235 VSS.n65 8.84261
R1248 VSS.n2180 VSS.n170 8.84261
R1249 VSS.n703 VSS.n587 8.41029
R1250 VSS.n1848 VSS.n1847 8.16291
R1251 VSS.n1903 VSS.n1902 8.04205
R1252 VSS.n1821 VSS.n233 8.03936
R1253 VSS.n570 VSS.n567 7.92155
R1254 VSS.n516 VSS.n513 7.92155
R1255 VSS.n463 VSS.n443 7.92155
R1256 VSS.n421 VSS.n368 7.92155
R1257 VSS.n10 VSS.n7 7.92155
R1258 VSS.n2291 VSS.n49 7.92155
R1259 VSS.n80 VSS.n61 7.92155
R1260 VSS.n2101 VSS.t1 7.84851
R1261 VSS.n673 VSS.n621 7.82945
R1262 VSS.n1206 VSS.n588 7.82945
R1263 VSS.n1334 VSS.n534 7.82945
R1264 VSS.n1495 VSS.n481 7.82945
R1265 VSS.n381 VSS.n328 7.82945
R1266 VSS.n2342 VSS.n28 7.82945
R1267 VSS.n1836 VSS.n248 7.82945
R1268 VSS.n2176 VSS.n170 7.82945
R1269 VSS.n121 VSS.n65 7.82945
R1270 VSS.n2049 VSS.n2030 6.44787
R1271 VSS.n1727 VSS.n283 6.44787
R1272 VSS.n1644 VSS.n307 6.44787
R1273 VSS.n875 VSS.n830 6.44787
R1274 VSS.n812 VSS.n720 6.44787
R1275 VSS.n1026 VSS.n994 6.44787
R1276 VSS.n1759 VSS.n217 6.44787
R1277 VSS.n1132 VSS.n604 6.28069
R1278 VSS.n1260 VSS.n550 6.28069
R1279 VSS.n1388 VSS.n497 6.28069
R1280 VSS.n1449 VSS.n1448 6.28069
R1281 VSS.n1591 VSS.n1590 6.28069
R1282 VSS.n2296 VSS.n2295 6.28069
R1283 VSS.n766 VSS.n703 6.05199
R1284 VSS.n1907 VSS.n1906 5.99128
R1285 VSS.n1951 VSS.n223 5.99128
R1286 VSS.n1948 VSS.n1947 5.99128
R1287 VSS.n1913 VSS.n229 5.99128
R1288 VSS.n1941 VSS.n1914 5.99128
R1289 VSS.n1940 VSS.n1915 5.99128
R1290 VSS.n1923 VSS.n1922 5.99128
R1291 VSS.n1934 VSS.n1933 5.99128
R1292 VSS.n1927 VSS.n1924 5.99128
R1293 VSS.n1926 VSS.n62 5.99128
R1294 VSS.n2237 VSS.n2236 5.99128
R1295 VSS.n2230 VSS.n126 5.99128
R1296 VSS.n2229 VSS.n127 5.99128
R1297 VSS.n2226 VSS.n2225 5.99128
R1298 VSS.n134 VSS.n130 5.99128
R1299 VSS.n2219 VSS.n135 5.99128
R1300 VSS.n2218 VSS.n136 5.99128
R1301 VSS.n1132 VSS.n1131 5.58327
R1302 VSS.n1260 VSS.n1259 5.58327
R1303 VSS.n1388 VSS.n1387 5.58327
R1304 VSS.n1448 VSS.n436 5.58327
R1305 VSS.n1590 VSS.n341 5.58327
R1306 VSS.n2295 VSS.n43 5.58327
R1307 VSS.n2209 VSS.n2208 5.54027
R1308 VSS.n2102 VSS.n2101 5.54027
R1309 VSS.n2202 VSS.n150 5.54027
R1310 VSS.n2201 VSS.n151 5.54027
R1311 VSS.n2127 VSS.n158 5.54027
R1312 VSS.n2195 VSS.n2194 5.54027
R1313 VSS.n2077 VSS.n159 5.54027
R1314 VSS.n2188 VSS.n165 5.54027
R1315 VSS.n2187 VSS.n166 5.54027
R1316 VSS.n2182 VSS.n2181 5.54027
R1317 VSS.n1003 VSS.n1002 5.2005
R1318 VSS.n1005 VSS.n1004 5.2005
R1319 VSS.n1007 VSS.n1006 5.2005
R1320 VSS.n1009 VSS.n1008 5.2005
R1321 VSS.n1011 VSS.n1010 5.2005
R1322 VSS.n1013 VSS.n1012 5.2005
R1323 VSS.n1015 VSS.n1014 5.2005
R1324 VSS.n1017 VSS.n1016 5.2005
R1325 VSS.n1019 VSS.n1018 5.2005
R1326 VSS.n1021 VSS.n1020 5.2005
R1327 VSS.n1023 VSS.n1022 5.2005
R1328 VSS.n1024 VSS.n995 5.2005
R1329 VSS.n1026 VSS.n1025 5.2005
R1330 VSS.n1027 VSS.n1026 5.2005
R1331 VSS.n789 VSS.n788 5.2005
R1332 VSS.n788 VSS.n787 5.2005
R1333 VSS.n790 VSS.n780 5.2005
R1334 VSS.n780 VSS.n779 5.2005
R1335 VSS.n792 VSS.n791 5.2005
R1336 VSS.n793 VSS.n792 5.2005
R1337 VSS.n777 VSS.n776 5.2005
R1338 VSS.n794 VSS.n777 5.2005
R1339 VSS.n797 VSS.n796 5.2005
R1340 VSS.n796 VSS.n795 5.2005
R1341 VSS.n798 VSS.n775 5.2005
R1342 VSS.n775 VSS.n774 5.2005
R1343 VSS.n800 VSS.n799 5.2005
R1344 VSS.n801 VSS.n800 5.2005
R1345 VSS.n773 VSS.n772 5.2005
R1346 VSS.n802 VSS.n773 5.2005
R1347 VSS.n805 VSS.n804 5.2005
R1348 VSS.n804 VSS.n803 5.2005
R1349 VSS.n806 VSS.n771 5.2005
R1350 VSS.n771 VSS.n770 5.2005
R1351 VSS.n808 VSS.n807 5.2005
R1352 VSS.n809 VSS.n808 5.2005
R1353 VSS.n769 VSS.n768 5.2005
R1354 VSS.n810 VSS.n769 5.2005
R1355 VSS.n813 VSS.n812 5.2005
R1356 VSS.n812 VSS.n811 5.2005
R1357 VSS.n852 VSS.n851 5.2005
R1358 VSS.n851 VSS.n850 5.2005
R1359 VSS.n853 VSS.n843 5.2005
R1360 VSS.n843 VSS.n842 5.2005
R1361 VSS.n855 VSS.n854 5.2005
R1362 VSS.n856 VSS.n855 5.2005
R1363 VSS.n841 VSS.n840 5.2005
R1364 VSS.n857 VSS.n841 5.2005
R1365 VSS.n860 VSS.n859 5.2005
R1366 VSS.n859 VSS.n858 5.2005
R1367 VSS.n861 VSS.n839 5.2005
R1368 VSS.n839 VSS.n838 5.2005
R1369 VSS.n863 VSS.n862 5.2005
R1370 VSS.n864 VSS.n863 5.2005
R1371 VSS.n837 VSS.n836 5.2005
R1372 VSS.n865 VSS.n837 5.2005
R1373 VSS.n868 VSS.n867 5.2005
R1374 VSS.n867 VSS.n866 5.2005
R1375 VSS.n869 VSS.n835 5.2005
R1376 VSS.n835 VSS.n834 5.2005
R1377 VSS.n871 VSS.n870 5.2005
R1378 VSS.n872 VSS.n871 5.2005
R1379 VSS.n833 VSS.n832 5.2005
R1380 VSS.n873 VSS.n833 5.2005
R1381 VSS.n876 VSS.n875 5.2005
R1382 VSS.n875 VSS.n874 5.2005
R1383 VSS.n1619 VSS.n1618 5.2005
R1384 VSS.n1620 VSS.n1619 5.2005
R1385 VSS.n322 VSS.n321 5.2005
R1386 VSS.n1621 VSS.n322 5.2005
R1387 VSS.n1624 VSS.n1623 5.2005
R1388 VSS.n1623 VSS.n1622 5.2005
R1389 VSS.n1625 VSS.n320 5.2005
R1390 VSS.n320 VSS.n319 5.2005
R1391 VSS.n1627 VSS.n1626 5.2005
R1392 VSS.n1628 VSS.n1627 5.2005
R1393 VSS.n317 VSS.n316 5.2005
R1394 VSS.n1630 VSS.n317 5.2005
R1395 VSS.n1633 VSS.n1632 5.2005
R1396 VSS.n1632 VSS.n1631 5.2005
R1397 VSS.n1634 VSS.n315 5.2005
R1398 VSS.n315 VSS.n314 5.2005
R1399 VSS.n1636 VSS.n1635 5.2005
R1400 VSS.n1637 VSS.n1636 5.2005
R1401 VSS.n313 VSS.n312 5.2005
R1402 VSS.n1638 VSS.n313 5.2005
R1403 VSS.n1641 VSS.n1640 5.2005
R1404 VSS.n1640 VSS.n1639 5.2005
R1405 VSS.n1642 VSS.n308 5.2005
R1406 VSS.n308 VSS.n306 5.2005
R1407 VSS.n1644 VSS.n1643 5.2005
R1408 VSS.n1645 VSS.n1644 5.2005
R1409 VSS.n1704 VSS.n1703 5.2005
R1410 VSS.n1703 VSS.n1702 5.2005
R1411 VSS.n1705 VSS.n1694 5.2005
R1412 VSS.n1694 VSS.n1693 5.2005
R1413 VSS.n1707 VSS.n1706 5.2005
R1414 VSS.n1708 VSS.n1707 5.2005
R1415 VSS.n1695 VSS.n1691 5.2005
R1416 VSS.n1709 VSS.n1691 5.2005
R1417 VSS.n1711 VSS.n1692 5.2005
R1418 VSS.n1711 VSS.n1710 5.2005
R1419 VSS.n1712 VSS.n1690 5.2005
R1420 VSS.n1713 VSS.n1712 5.2005
R1421 VSS.n1716 VSS.n1715 5.2005
R1422 VSS.n1715 VSS.n1714 5.2005
R1423 VSS.n1717 VSS.n1689 5.2005
R1424 VSS.n1689 VSS.n1688 5.2005
R1425 VSS.n1719 VSS.n1718 5.2005
R1426 VSS.n1720 VSS.n1719 5.2005
R1427 VSS.n1687 VSS.n1686 5.2005
R1428 VSS.n1721 VSS.n1687 5.2005
R1429 VSS.n1724 VSS.n1723 5.2005
R1430 VSS.n1723 VSS.n1722 5.2005
R1431 VSS.n1725 VSS.n284 5.2005
R1432 VSS.n284 VSS.n282 5.2005
R1433 VSS.n1727 VSS.n1726 5.2005
R1434 VSS.n1728 VSS.n1727 5.2005
R1435 VSS.n10 VSS.n4 5.2005
R1436 VSS.n2349 VSS.n2348 5.2005
R1437 VSS.n2351 VSS.n2350 5.2005
R1438 VSS.n2352 VSS.n14 5.2005
R1439 VSS.n2354 VSS.n2353 5.2005
R1440 VSS.n2355 VSS.n2354 5.2005
R1441 VSS.n422 VSS.n421 5.2005
R1442 VSS.n419 VSS.n370 5.2005
R1443 VSS.n418 VSS.n417 5.2005
R1444 VSS.n416 VSS.n415 5.2005
R1445 VSS.n414 VSS.n372 5.2005
R1446 VSS.n414 VSS.n367 5.2005
R1447 VSS.n463 VSS.n440 5.2005
R1448 VSS.n1502 VSS.n1501 5.2005
R1449 VSS.n1504 VSS.n1503 5.2005
R1450 VSS.n1505 VSS.n467 5.2005
R1451 VSS.n1507 VSS.n1506 5.2005
R1452 VSS.n1508 VSS.n1507 5.2005
R1453 VSS.n516 VSS.n509 5.2005
R1454 VSS.n1341 VSS.n1340 5.2005
R1455 VSS.n1343 VSS.n1342 5.2005
R1456 VSS.n1344 VSS.n520 5.2005
R1457 VSS.n1346 VSS.n1345 5.2005
R1458 VSS.n1347 VSS.n1346 5.2005
R1459 VSS.n570 VSS.n563 5.2005
R1460 VSS.n1213 VSS.n1212 5.2005
R1461 VSS.n1215 VSS.n1214 5.2005
R1462 VSS.n1216 VSS.n574 5.2005
R1463 VSS.n1218 VSS.n1217 5.2005
R1464 VSS.n1219 VSS.n1218 5.2005
R1465 VSS.n641 VSS.n640 5.2005
R1466 VSS.n639 VSS.n638 5.2005
R1467 VSS.n637 VSS.n633 5.2005
R1468 VSS.n635 VSS.n634 5.2005
R1469 VSS.n617 VSS.n616 5.2005
R1470 VSS.n618 VSS.n617 5.2005
R1471 VSS.n591 VSS.n590 5.2005
R1472 VSS.n997 VSS.n996 5.2005
R1473 VSS.n999 VSS.n998 5.2005
R1474 VSS.n1001 VSS.n1000 5.2005
R1475 VSS.n537 VSS.n536 5.2005
R1476 VSS.n782 VSS.n781 5.2005
R1477 VSS.n784 VSS.n783 5.2005
R1478 VSS.n786 VSS.n785 5.2005
R1479 VSS.n484 VSS.n483 5.2005
R1480 VSS.n845 VSS.n844 5.2005
R1481 VSS.n847 VSS.n846 5.2005
R1482 VSS.n849 VSS.n848 5.2005
R1483 VSS.n1612 VSS.n1611 5.2005
R1484 VSS.n1614 VSS.n325 5.2005
R1485 VSS.n1616 VSS.n1615 5.2005
R1486 VSS.n1617 VSS.n324 5.2005
R1487 VSS.n31 VSS.n30 5.2005
R1488 VSS.n1697 VSS.n1696 5.2005
R1489 VSS.n1699 VSS.n1698 5.2005
R1490 VSS.n1701 VSS.n1700 5.2005
R1491 VSS.n674 VSS.n673 5.2005
R1492 VSS.n671 VSS.n623 5.2005
R1493 VSS.n670 VSS.n669 5.2005
R1494 VSS.n668 VSS.n667 5.2005
R1495 VSS.n666 VSS.n625 5.2005
R1496 VSS.n664 VSS.n663 5.2005
R1497 VSS.n662 VSS.n626 5.2005
R1498 VSS.n661 VSS.n660 5.2005
R1499 VSS.n658 VSS.n627 5.2005
R1500 VSS.n656 VSS.n655 5.2005
R1501 VSS.n654 VSS.n628 5.2005
R1502 VSS.n653 VSS.n652 5.2005
R1503 VSS.n650 VSS.n629 5.2005
R1504 VSS.n648 VSS.n647 5.2005
R1505 VSS.n646 VSS.n630 5.2005
R1506 VSS.n645 VSS.n644 5.2005
R1507 VSS.n642 VSS.n631 5.2005
R1508 VSS.n642 VSS.n619 5.2005
R1509 VSS.n1211 VSS.n573 5.2005
R1510 VSS.n1210 VSS.n1209 5.2005
R1511 VSS.n576 VSS.n575 5.2005
R1512 VSS.n1181 VSS.n1180 5.2005
R1513 VSS.n1183 VSS.n1182 5.2005
R1514 VSS.n1185 VSS.n1184 5.2005
R1515 VSS.n1187 VSS.n1186 5.2005
R1516 VSS.n1189 VSS.n1188 5.2005
R1517 VSS.n1191 VSS.n1190 5.2005
R1518 VSS.n1193 VSS.n1192 5.2005
R1519 VSS.n1195 VSS.n1194 5.2005
R1520 VSS.n1197 VSS.n1196 5.2005
R1521 VSS.n1199 VSS.n1198 5.2005
R1522 VSS.n1201 VSS.n1200 5.2005
R1523 VSS.n1203 VSS.n1202 5.2005
R1524 VSS.n1204 VSS.n589 5.2005
R1525 VSS.n1206 VSS.n1205 5.2005
R1526 VSS.n1207 VSS.n1206 5.2005
R1527 VSS.n1339 VSS.n519 5.2005
R1528 VSS.n1338 VSS.n1337 5.2005
R1529 VSS.n522 VSS.n521 5.2005
R1530 VSS.n1309 VSS.n1308 5.2005
R1531 VSS.n1311 VSS.n1310 5.2005
R1532 VSS.n1313 VSS.n1312 5.2005
R1533 VSS.n1315 VSS.n1314 5.2005
R1534 VSS.n1317 VSS.n1316 5.2005
R1535 VSS.n1319 VSS.n1318 5.2005
R1536 VSS.n1321 VSS.n1320 5.2005
R1537 VSS.n1323 VSS.n1322 5.2005
R1538 VSS.n1325 VSS.n1324 5.2005
R1539 VSS.n1327 VSS.n1326 5.2005
R1540 VSS.n1329 VSS.n1328 5.2005
R1541 VSS.n1331 VSS.n1330 5.2005
R1542 VSS.n1332 VSS.n535 5.2005
R1543 VSS.n1334 VSS.n1333 5.2005
R1544 VSS.n1335 VSS.n1334 5.2005
R1545 VSS.n1500 VSS.n466 5.2005
R1546 VSS.n1499 VSS.n1498 5.2005
R1547 VSS.n469 VSS.n468 5.2005
R1548 VSS.n1470 VSS.n1469 5.2005
R1549 VSS.n1472 VSS.n1471 5.2005
R1550 VSS.n1474 VSS.n1473 5.2005
R1551 VSS.n1476 VSS.n1475 5.2005
R1552 VSS.n1478 VSS.n1477 5.2005
R1553 VSS.n1480 VSS.n1479 5.2005
R1554 VSS.n1482 VSS.n1481 5.2005
R1555 VSS.n1484 VSS.n1483 5.2005
R1556 VSS.n1486 VSS.n1485 5.2005
R1557 VSS.n1488 VSS.n1487 5.2005
R1558 VSS.n1490 VSS.n1489 5.2005
R1559 VSS.n1492 VSS.n1491 5.2005
R1560 VSS.n1493 VSS.n482 5.2005
R1561 VSS.n1495 VSS.n1494 5.2005
R1562 VSS.n1496 VSS.n1495 5.2005
R1563 VSS.n413 VSS.n373 5.2005
R1564 VSS.n411 VSS.n410 5.2005
R1565 VSS.n409 VSS.n374 5.2005
R1566 VSS.n408 VSS.n407 5.2005
R1567 VSS.n405 VSS.n375 5.2005
R1568 VSS.n403 VSS.n402 5.2005
R1569 VSS.n401 VSS.n376 5.2005
R1570 VSS.n400 VSS.n399 5.2005
R1571 VSS.n397 VSS.n377 5.2005
R1572 VSS.n395 VSS.n394 5.2005
R1573 VSS.n393 VSS.n378 5.2005
R1574 VSS.n392 VSS.n391 5.2005
R1575 VSS.n389 VSS.n379 5.2005
R1576 VSS.n387 VSS.n386 5.2005
R1577 VSS.n385 VSS.n380 5.2005
R1578 VSS.n384 VSS.n383 5.2005
R1579 VSS.n381 VSS.n329 5.2005
R1580 VSS.n381 VSS.n327 5.2005
R1581 VSS.n2347 VSS.n13 5.2005
R1582 VSS.n2346 VSS.n2345 5.2005
R1583 VSS.n16 VSS.n15 5.2005
R1584 VSS.n2317 VSS.n2316 5.2005
R1585 VSS.n2319 VSS.n2318 5.2005
R1586 VSS.n2321 VSS.n2320 5.2005
R1587 VSS.n2323 VSS.n2322 5.2005
R1588 VSS.n2325 VSS.n2324 5.2005
R1589 VSS.n2327 VSS.n2326 5.2005
R1590 VSS.n2329 VSS.n2328 5.2005
R1591 VSS.n2331 VSS.n2330 5.2005
R1592 VSS.n2333 VSS.n2332 5.2005
R1593 VSS.n2335 VSS.n2334 5.2005
R1594 VSS.n2337 VSS.n2336 5.2005
R1595 VSS.n2339 VSS.n2338 5.2005
R1596 VSS.n2340 VSS.n29 5.2005
R1597 VSS.n2342 VSS.n2341 5.2005
R1598 VSS.n2343 VSS.n2342 5.2005
R1599 VSS.n2015 VSS.n2014 5.2005
R1600 VSS.n2014 VSS.n2013 5.2005
R1601 VSS.n2016 VSS.n1992 5.2005
R1602 VSS.n1992 VSS.n1991 5.2005
R1603 VSS.n2018 VSS.n2017 5.2005
R1604 VSS.n2019 VSS.n2018 5.2005
R1605 VSS.n1990 VSS.n1989 5.2005
R1606 VSS.n2020 VSS.n1990 5.2005
R1607 VSS.n2023 VSS.n2022 5.2005
R1608 VSS.n2022 VSS.n2021 5.2005
R1609 VSS.n2024 VSS.n1987 5.2005
R1610 VSS.n1987 VSS.n1986 5.2005
R1611 VSS.n2026 VSS.n2025 5.2005
R1612 VSS.n2027 VSS.n2026 5.2005
R1613 VSS.n1988 VSS.n1984 5.2005
R1614 VSS.n2028 VSS.n1984 5.2005
R1615 VSS.n2030 VSS.n1985 5.2005
R1616 VSS.n2030 VSS.n2029 5.2005
R1617 VSS.n1997 VSS.n123 5.2005
R1618 VSS.n2000 VSS.n1999 5.2005
R1619 VSS.n2002 VSS.n2001 5.2005
R1620 VSS.n2004 VSS.n1995 5.2005
R1621 VSS.n2006 VSS.n2005 5.2005
R1622 VSS.n2007 VSS.n1994 5.2005
R1623 VSS.n2009 VSS.n2008 5.2005
R1624 VSS.n2011 VSS.n1993 5.2005
R1625 VSS.n2096 VSS.n2095 5.2005
R1626 VSS.n2094 VSS.n2093 5.2005
R1627 VSS.n2092 VSS.n178 5.2005
R1628 VSS.n2086 VSS.n179 5.2005
R1629 VSS.n2088 VSS.n2087 5.2005
R1630 VSS.n2085 VSS.n181 5.2005
R1631 VSS.n2100 VSS.n2099 5.2005
R1632 VSS.n2097 VSS.n176 5.2005
R1633 VSS.n2121 VSS.n2120 5.2005
R1634 VSS.n2118 VSS.n171 5.2005
R1635 VSS.n2117 VSS.n172 5.2005
R1636 VSS.n2115 VSS.n2114 5.2005
R1637 VSS.n2113 VSS.n173 5.2005
R1638 VSS.n2112 VSS.n2111 5.2005
R1639 VSS.n2109 VSS.n174 5.2005
R1640 VSS.n2107 VSS.n2106 5.2005
R1641 VSS.n2105 VSS.n175 5.2005
R1642 VSS.n175 VSS.n169 5.2005
R1643 VSS.n723 VSS.n722 5.2005
R1644 VSS.n739 VSS.n723 5.2005
R1645 VSS.n737 VSS.n736 5.2005
R1646 VSS.n738 VSS.n737 5.2005
R1647 VSS.n735 VSS.n725 5.2005
R1648 VSS.n725 VSS.n724 5.2005
R1649 VSS.n734 VSS.n733 5.2005
R1650 VSS.n733 VSS.n732 5.2005
R1651 VSS.n727 VSS.n726 5.2005
R1652 VSS.n731 VSS.n727 5.2005
R1653 VSS.n729 VSS.n728 5.2005
R1654 VSS.n730 VSS.n729 5.2005
R1655 VSS.n683 VSS.n682 5.2005
R1656 VSS.n684 VSS.n683 5.2005
R1657 VSS.n1048 VSS.n1047 5.2005
R1658 VSS.n1047 VSS.n1046 5.2005
R1659 VSS.n1049 VSS.n681 5.2005
R1660 VSS.n681 VSS.n680 5.2005
R1661 VSS.n1051 VSS.n1050 5.2005
R1662 VSS.n1052 VSS.n1051 5.2005
R1663 VSS.n679 VSS.n678 5.2005
R1664 VSS.n1053 VSS.n679 5.2005
R1665 VSS.n1057 VSS.n1056 5.2005
R1666 VSS.n1056 VSS.n1055 5.2005
R1667 VSS.n1058 VSS.n677 5.2005
R1668 VSS.n1054 VSS.n677 5.2005
R1669 VSS.n1060 VSS.n1059 5.2005
R1670 VSS.n1062 VSS.n676 5.2005
R1671 VSS.n1063 VSS.n675 5.2005
R1672 VSS.n1066 VSS.n1065 5.2005
R1673 VSS.n2084 VSS.n185 5.2005
R1674 VSS.n2080 VSS.n185 5.2005
R1675 VSS.n2083 VSS.n2082 5.2005
R1676 VSS.n2082 VSS.n2081 5.2005
R1677 VSS.n187 VSS.n186 5.2005
R1678 VSS.n2079 VSS.n187 5.2005
R1679 VSS.n2075 VSS.n2074 5.2005
R1680 VSS.n2076 VSS.n2075 5.2005
R1681 VSS.n2073 VSS.n189 5.2005
R1682 VSS.n189 VSS.n188 5.2005
R1683 VSS.n2072 VSS.n2071 5.2005
R1684 VSS.n2071 VSS.n2070 5.2005
R1685 VSS.n191 VSS.n190 5.2005
R1686 VSS.n2069 VSS.n191 5.2005
R1687 VSS.n2067 VSS.n2066 5.2005
R1688 VSS.n2068 VSS.n2067 5.2005
R1689 VSS.n2065 VSS.n193 5.2005
R1690 VSS.n193 VSS.n192 5.2005
R1691 VSS.n2064 VSS.n2063 5.2005
R1692 VSS.n195 VSS.n194 5.2005
R1693 VSS.n2034 VSS.n2032 5.2005
R1694 VSS.n2035 VSS.n2031 5.2005
R1695 VSS.n2035 VSS.n196 5.2005
R1696 VSS.n2037 VSS.n2036 5.2005
R1697 VSS.n2039 VSS.n2038 5.2005
R1698 VSS.n2041 VSS.n2040 5.2005
R1699 VSS.n2043 VSS.n2042 5.2005
R1700 VSS.n2045 VSS.n2044 5.2005
R1701 VSS.n2048 VSS.n2047 5.2005
R1702 VSS.n2051 VSS.n2050 5.2005
R1703 VSS.n2054 VSS.n2053 5.2005
R1704 VSS.n2056 VSS.n2055 5.2005
R1705 VSS.n2057 VSS.n214 5.2005
R1706 VSS.n2059 VSS.n2058 5.2005
R1707 VSS.n2060 VSS.n2059 5.2005
R1708 VSS.n215 VSS.n213 5.2005
R1709 VSS.n1959 VSS.n1958 5.2005
R1710 VSS.n1961 VSS.n1960 5.2005
R1711 VSS.n1963 VSS.n1955 5.2005
R1712 VSS.n1965 VSS.n1964 5.2005
R1713 VSS.n1966 VSS.n1954 5.2005
R1714 VSS.n1968 VSS.n1967 5.2005
R1715 VSS.n1970 VSS.n221 5.2005
R1716 VSS.n1972 VSS.n1971 5.2005
R1717 VSS.n1973 VSS.n220 5.2005
R1718 VSS.n1975 VSS.n1974 5.2005
R1719 VSS.n1977 VSS.n219 5.2005
R1720 VSS.n1978 VSS.n216 5.2005
R1721 VSS.n1981 VSS.n1980 5.2005
R1722 VSS.n1756 VSS.n1755 5.2005
R1723 VSS.n1753 VSS.n1752 5.2005
R1724 VSS.n1751 VSS.n267 5.2005
R1725 VSS.n1750 VSS.n1749 5.2005
R1726 VSS.n1747 VSS.n268 5.2005
R1727 VSS.n1745 VSS.n1744 5.2005
R1728 VSS.n1743 VSS.n269 5.2005
R1729 VSS.n1742 VSS.n1741 5.2005
R1730 VSS.n1739 VSS.n270 5.2005
R1731 VSS.n1734 VSS.n271 5.2005
R1732 VSS.n1736 VSS.n1735 5.2005
R1733 VSS.n1737 VSS.n1736 5.2005
R1734 VSS.n1733 VSS.n272 5.2005
R1735 VSS.n1732 VSS.n1731 5.2005
R1736 VSS.n274 VSS.n273 5.2005
R1737 VSS.n1675 VSS.n1674 5.2005
R1738 VSS.n1677 VSS.n1676 5.2005
R1739 VSS.n1679 VSS.n1678 5.2005
R1740 VSS.n1681 VSS.n1680 5.2005
R1741 VSS.n1684 VSS.n1683 5.2005
R1742 VSS.n1673 VSS.n1672 5.2005
R1743 VSS.n1670 VSS.n1669 5.2005
R1744 VSS.n1668 VSS.n1667 5.2005
R1745 VSS.n1666 VSS.n1665 5.2005
R1746 VSS.n1664 VSS.n1663 5.2005
R1747 VSS.n1662 VSS.n1661 5.2005
R1748 VSS.n1660 VSS.n1659 5.2005
R1749 VSS.n1658 VSS.n1657 5.2005
R1750 VSS.n1656 VSS.n286 5.2005
R1751 VSS.n1651 VSS.n287 5.2005
R1752 VSS.n1653 VSS.n1652 5.2005
R1753 VSS.n1654 VSS.n1653 5.2005
R1754 VSS.n1650 VSS.n288 5.2005
R1755 VSS.n1649 VSS.n1648 5.2005
R1756 VSS.n290 VSS.n289 5.2005
R1757 VSS.n304 VSS.n303 5.2005
R1758 VSS.n302 VSS.n297 5.2005
R1759 VSS.n301 VSS.n300 5.2005
R1760 VSS.n299 VSS.n298 5.2005
R1761 VSS.n310 VSS.n309 5.2005
R1762 VSS.n888 VSS.n887 5.2005
R1763 VSS.n891 VSS.n890 5.2005
R1764 VSS.n893 VSS.n892 5.2005
R1765 VSS.n895 VSS.n894 5.2005
R1766 VSS.n897 VSS.n896 5.2005
R1767 VSS.n899 VSS.n898 5.2005
R1768 VSS.n901 VSS.n900 5.2005
R1769 VSS.n902 VSS.n885 5.2005
R1770 VSS.n904 VSS.n903 5.2005
R1771 VSS.n886 VSS.n884 5.2005
R1772 VSS.n907 VSS.n882 5.2005
R1773 VSS.n907 VSS.n906 5.2005
R1774 VSS.n909 VSS.n908 5.2005
R1775 VSS.n910 VSS.n881 5.2005
R1776 VSS.n912 VSS.n911 5.2005
R1777 VSS.n914 VSS.n879 5.2005
R1778 VSS.n916 VSS.n915 5.2005
R1779 VSS.n917 VSS.n878 5.2005
R1780 VSS.n919 VSS.n918 5.2005
R1781 VSS.n922 VSS.n921 5.2005
R1782 VSS.n925 VSS.n924 5.2005
R1783 VSS.n927 VSS.n828 5.2005
R1784 VSS.n929 VSS.n928 5.2005
R1785 VSS.n930 VSS.n827 5.2005
R1786 VSS.n932 VSS.n931 5.2005
R1787 VSS.n934 VSS.n824 5.2005
R1788 VSS.n936 VSS.n935 5.2005
R1789 VSS.n937 VSS.n822 5.2005
R1790 VSS.n939 VSS.n938 5.2005
R1791 VSS.n823 VSS.n821 5.2005
R1792 VSS.n942 VSS.n819 5.2005
R1793 VSS.n942 VSS.n941 5.2005
R1794 VSS.n944 VSS.n943 5.2005
R1795 VSS.n945 VSS.n818 5.2005
R1796 VSS.n947 VSS.n946 5.2005
R1797 VSS.n949 VSS.n816 5.2005
R1798 VSS.n951 VSS.n950 5.2005
R1799 VSS.n952 VSS.n815 5.2005
R1800 VSS.n954 VSS.n953 5.2005
R1801 VSS.n957 VSS.n956 5.2005
R1802 VSS.n960 VSS.n959 5.2005
R1803 VSS.n962 VSS.n718 5.2005
R1804 VSS.n964 VSS.n963 5.2005
R1805 VSS.n965 VSS.n717 5.2005
R1806 VSS.n967 VSS.n966 5.2005
R1807 VSS.n969 VSS.n714 5.2005
R1808 VSS.n971 VSS.n970 5.2005
R1809 VSS.n972 VSS.n713 5.2005
R1810 VSS.n974 VSS.n973 5.2005
R1811 VSS.n712 VSS.n711 5.2005
R1812 VSS.n978 VSS.n977 5.2005
R1813 VSS.n977 VSS.n976 5.2005
R1814 VSS.n979 VSS.n710 5.2005
R1815 VSS.n710 VSS.n709 5.2005
R1816 VSS.n981 VSS.n980 5.2005
R1817 VSS.n982 VSS.n981 5.2005
R1818 VSS.n708 VSS.n707 5.2005
R1819 VSS.n983 VSS.n708 5.2005
R1820 VSS.n986 VSS.n985 5.2005
R1821 VSS.n985 VSS.n984 5.2005
R1822 VSS.n987 VSS.n705 5.2005
R1823 VSS.n705 VSS.n704 5.2005
R1824 VSS.n989 VSS.n988 5.2005
R1825 VSS.n990 VSS.n989 5.2005
R1826 VSS.n706 VSS.n702 5.2005
R1827 VSS.n991 VSS.n702 5.2005
R1828 VSS.n993 VSS.n694 5.2005
R1829 VSS.n993 VSS.n992 5.2005
R1830 VSS.n695 VSS.n694 5.2005
R1831 VSS.n1028 VSS.n695 5.2005
R1832 VSS.n1031 VSS.n1030 5.2005
R1833 VSS.n1030 VSS.n1029 5.2005
R1834 VSS.n1032 VSS.n693 5.2005
R1835 VSS.n693 VSS.n692 5.2005
R1836 VSS.n1034 VSS.n1033 5.2005
R1837 VSS.n1035 VSS.n1034 5.2005
R1838 VSS.n691 VSS.n690 5.2005
R1839 VSS.n1036 VSS.n691 5.2005
R1840 VSS.n1039 VSS.n1038 5.2005
R1841 VSS.n1038 VSS.n1037 5.2005
R1842 VSS.n1040 VSS.n688 5.2005
R1843 VSS.n688 VSS.n686 5.2005
R1844 VSS.n1042 VSS.n1041 5.2005
R1845 VSS.n1043 VSS.n1042 5.2005
R1846 VSS.n689 VSS.n687 5.2005
R1847 VSS.n687 VSS.n685 5.2005
R1848 VSS.n749 VSS.n748 5.2005
R1849 VSS.n748 VSS.n747 5.2005
R1850 VSS.n750 VSS.n745 5.2005
R1851 VSS.n746 VSS.n745 5.2005
R1852 VSS.n752 VSS.n751 5.2005
R1853 VSS.n754 VSS.n743 5.2005
R1854 VSS.n756 VSS.n755 5.2005
R1855 VSS.n757 VSS.n742 5.2005
R1856 VSS.n759 VSS.n758 5.2005
R1857 VSS.n761 VSS.n741 5.2005
R1858 VSS.n762 VSS.n721 5.2005
R1859 VSS.n765 VSS.n764 5.2005
R1860 VSS.n1793 VSS.n1792 5.2005
R1861 VSS.n1792 VSS.n1791 5.2005
R1862 VSS.n250 VSS.n249 5.2005
R1863 VSS.n1790 VSS.n250 5.2005
R1864 VSS.n1788 VSS.n1787 5.2005
R1865 VSS.n1789 VSS.n1788 5.2005
R1866 VSS.n1786 VSS.n252 5.2005
R1867 VSS.n252 VSS.n251 5.2005
R1868 VSS.n1785 VSS.n1784 5.2005
R1869 VSS.n1784 VSS.n1783 5.2005
R1870 VSS.n254 VSS.n253 5.2005
R1871 VSS.n1782 VSS.n254 5.2005
R1872 VSS.n1780 VSS.n1779 5.2005
R1873 VSS.n1781 VSS.n1780 5.2005
R1874 VSS.n1778 VSS.n256 5.2005
R1875 VSS.n256 VSS.n255 5.2005
R1876 VSS.n1777 VSS.n1776 5.2005
R1877 VSS.n1776 VSS.n1775 5.2005
R1878 VSS.n258 VSS.n257 5.2005
R1879 VSS.n1773 VSS.n258 5.2005
R1880 VSS.n1771 VSS.n1770 5.2005
R1881 VSS.n1772 VSS.n1771 5.2005
R1882 VSS.n1769 VSS.n261 5.2005
R1883 VSS.n261 VSS.n260 5.2005
R1884 VSS.n1768 VSS.n1767 5.2005
R1885 VSS.n1767 VSS.n1766 5.2005
R1886 VSS.n263 VSS.n262 5.2005
R1887 VSS.n1765 VSS.n263 5.2005
R1888 VSS.n1763 VSS.n1762 5.2005
R1889 VSS.n1764 VSS.n1763 5.2005
R1890 VSS.n1761 VSS.n265 5.2005
R1891 VSS.n265 VSS.n264 5.2005
R1892 VSS.n1760 VSS.n1759 5.2005
R1893 VSS.n1759 VSS.n1758 5.2005
R1894 VSS.n2291 VSS.n2290 5.2005
R1895 VSS.n2292 VSS.n2291 5.2005
R1896 VSS.n50 VSS.n48 5.2005
R1897 VSS.n48 VSS.n46 5.2005
R1898 VSS.n1861 VSS.n1860 5.2005
R1899 VSS.n1862 VSS.n1861 5.2005
R1900 VSS.n1865 VSS.n1864 5.2005
R1901 VSS.n1864 VSS.n1863 5.2005
R1902 VSS.n1866 VSS.n1859 5.2005
R1903 VSS.n1859 VSS.n1858 5.2005
R1904 VSS.n1868 VSS.n1867 5.2005
R1905 VSS.n1869 VSS.n1868 5.2005
R1906 VSS.n1857 VSS.n1856 5.2005
R1907 VSS.n1870 VSS.n1857 5.2005
R1908 VSS.n1873 VSS.n1872 5.2005
R1909 VSS.n1872 VSS.n1871 5.2005
R1910 VSS.n1874 VSS.n1855 5.2005
R1911 VSS.n1855 VSS.n1854 5.2005
R1912 VSS.n1876 VSS.n1875 5.2005
R1913 VSS.n1877 VSS.n1876 5.2005
R1914 VSS.n1853 VSS.n1852 5.2005
R1915 VSS.n1878 VSS.n1853 5.2005
R1916 VSS.n1881 VSS.n1880 5.2005
R1917 VSS.n1880 VSS.n1879 5.2005
R1918 VSS.n1882 VSS.n239 5.2005
R1919 VSS.n239 VSS.n237 5.2005
R1920 VSS.n1884 VSS.n1883 5.2005
R1921 VSS.n1885 VSS.n1884 5.2005
R1922 VSS.n1851 VSS.n238 5.2005
R1923 VSS.n238 VSS.n236 5.2005
R1924 VSS.n1850 VSS.n1849 5.2005
R1925 VSS.n1849 VSS.n1848 5.2005
R1926 VSS.n241 VSS.n240 5.2005
R1927 VSS.n1846 VSS.n241 5.2005
R1928 VSS.n1844 VSS.n1843 5.2005
R1929 VSS.n1845 VSS.n1844 5.2005
R1930 VSS.n1842 VSS.n244 5.2005
R1931 VSS.n244 VSS.n243 5.2005
R1932 VSS.n1841 VSS.n1840 5.2005
R1933 VSS.n1840 VSS.n1839 5.2005
R1934 VSS.n246 VSS.n245 5.2005
R1935 VSS.n1838 VSS.n246 5.2005
R1936 VSS.n1836 VSS.n1835 5.2005
R1937 VSS.n1837 VSS.n1836 5.2005
R1938 VSS.n2180 VSS.n2179 5.2005
R1939 VSS.n2181 VSS.n2180 5.2005
R1940 VSS.n164 VSS.n163 5.2005
R1941 VSS.n166 VSS.n164 5.2005
R1942 VSS.n2190 VSS.n2189 5.2005
R1943 VSS.n2189 VSS.n2188 5.2005
R1944 VSS.n2191 VSS.n161 5.2005
R1945 VSS.n2077 VSS.n161 5.2005
R1946 VSS.n2193 VSS.n2192 5.2005
R1947 VSS.n2194 VSS.n2193 5.2005
R1948 VSS.n162 VSS.n160 5.2005
R1949 VSS.n160 VSS.n158 5.2005
R1950 VSS.n149 VSS.n148 5.2005
R1951 VSS.n151 VSS.n149 5.2005
R1952 VSS.n2204 VSS.n2203 5.2005
R1953 VSS.n2203 VSS.n2202 5.2005
R1954 VSS.n2205 VSS.n146 5.2005
R1955 VSS.n2101 VSS.n146 5.2005
R1956 VSS.n2207 VSS.n2206 5.2005
R1957 VSS.n2208 VSS.n2207 5.2005
R1958 VSS.n147 VSS.n145 5.2005
R1959 VSS.n202 VSS.n201 5.2005
R1960 VSS.n204 VSS.n203 5.2005
R1961 VSS.n205 VSS.n204 5.2005
R1962 VSS.n133 VSS.n132 5.2005
R1963 VSS.n136 VSS.n133 5.2005
R1964 VSS.n2221 VSS.n2220 5.2005
R1965 VSS.n2220 VSS.n2219 5.2005
R1966 VSS.n2222 VSS.n131 5.2005
R1967 VSS.n134 VSS.n131 5.2005
R1968 VSS.n2224 VSS.n2223 5.2005
R1969 VSS.n2225 VSS.n2224 5.2005
R1970 VSS.n125 VSS.n124 5.2005
R1971 VSS.n127 VSS.n125 5.2005
R1972 VSS.n2232 VSS.n2231 5.2005
R1973 VSS.n2231 VSS.n2230 5.2005
R1974 VSS.n2235 VSS.n2234 5.2005
R1975 VSS.n2236 VSS.n2235 5.2005
R1976 VSS.n66 VSS.n64 5.2005
R1977 VSS.n64 VSS.n62 5.2005
R1978 VSS.n1930 VSS.n1928 5.2005
R1979 VSS.n1928 VSS.n1927 5.2005
R1980 VSS.n1932 VSS.n1931 5.2005
R1981 VSS.n1933 VSS.n1932 5.2005
R1982 VSS.n1929 VSS.n1925 5.2005
R1983 VSS.n1925 VSS.n1923 5.2005
R1984 VSS.n1912 VSS.n1911 5.2005
R1985 VSS.n1915 VSS.n1912 5.2005
R1986 VSS.n1943 VSS.n1942 5.2005
R1987 VSS.n1942 VSS.n1941 5.2005
R1988 VSS.n1944 VSS.n231 5.2005
R1989 VSS.n1913 VSS.n231 5.2005
R1990 VSS.n1946 VSS.n1945 5.2005
R1991 VSS.n1947 VSS.n1946 5.2005
R1992 VSS.n1910 VSS.n230 5.2005
R1993 VSS.n230 VSS.n223 5.2005
R1994 VSS.n1909 VSS.n1908 5.2005
R1995 VSS.n1908 VSS.n1907 5.2005
R1996 VSS.n233 VSS.n232 5.2005
R1997 VSS.n1822 VSS.n1819 5.2005
R1998 VSS.n1824 VSS.n1823 5.2005
R1999 VSS.n1825 VSS.n1818 5.2005
R2000 VSS.n1827 VSS.n1826 5.2005
R2001 VSS.n1829 VSS.n1817 5.2005
R2002 VSS.n1830 VSS.n1816 5.2005
R2003 VSS.n1833 VSS.n1832 5.2005
R2004 VSS.n1815 VSS.n1814 5.2005
R2005 VSS.n1812 VSS.n1794 5.2005
R2006 VSS.n1811 VSS.n1810 5.2005
R2007 VSS.n1809 VSS.n1808 5.2005
R2008 VSS.n1807 VSS.n1796 5.2005
R2009 VSS.n1805 VSS.n1804 5.2005
R2010 VSS.n1803 VSS.n1797 5.2005
R2011 VSS.n1802 VSS.n1801 5.2005
R2012 VSS.n1799 VSS.n1798 5.2005
R2013 VSS.n1799 VSS.n242 5.2005
R2014 VSS.n42 VSS.n41 5.2005
R2015 VSS.n44 VSS.n42 5.2005
R2016 VSS.n2298 VSS.n2297 5.2005
R2017 VSS.n2297 VSS.n2296 5.2005
R2018 VSS.n2299 VSS.n40 5.2005
R2019 VSS.n40 VSS.n39 5.2005
R2020 VSS.n2301 VSS.n2300 5.2005
R2021 VSS.n2302 VSS.n2301 5.2005
R2022 VSS.n38 VSS.n37 5.2005
R2023 VSS.n2303 VSS.n38 5.2005
R2024 VSS.n2306 VSS.n2305 5.2005
R2025 VSS.n2305 VSS.n2304 5.2005
R2026 VSS.n2307 VSS.n36 5.2005
R2027 VSS.n36 VSS.n35 5.2005
R2028 VSS.n2309 VSS.n2308 5.2005
R2029 VSS.n2310 VSS.n2309 5.2005
R2030 VSS.n34 VSS.n33 5.2005
R2031 VSS.n2311 VSS.n34 5.2005
R2032 VSS.n2314 VSS.n2313 5.2005
R2033 VSS.n2313 VSS.n2312 5.2005
R2034 VSS.n349 VSS.n32 5.2005
R2035 VSS.n349 VSS.n17 5.2005
R2036 VSS.n350 VSS.n348 5.2005
R2037 VSS.n1573 VSS.n350 5.2005
R2038 VSS.n1576 VSS.n1575 5.2005
R2039 VSS.n1575 VSS.n1574 5.2005
R2040 VSS.n1577 VSS.n347 5.2005
R2041 VSS.n347 VSS.n346 5.2005
R2042 VSS.n1579 VSS.n1578 5.2005
R2043 VSS.n1580 VSS.n1579 5.2005
R2044 VSS.n345 VSS.n344 5.2005
R2045 VSS.n1581 VSS.n345 5.2005
R2046 VSS.n1584 VSS.n1583 5.2005
R2047 VSS.n1583 VSS.n1582 5.2005
R2048 VSS.n1585 VSS.n343 5.2005
R2049 VSS.n343 VSS.n342 5.2005
R2050 VSS.n1587 VSS.n1586 5.2005
R2051 VSS.n1588 VSS.n1587 5.2005
R2052 VSS.n340 VSS.n339 5.2005
R2053 VSS.n1589 VSS.n340 5.2005
R2054 VSS.n1593 VSS.n1592 5.2005
R2055 VSS.n1592 VSS.n1591 5.2005
R2056 VSS.n1594 VSS.n338 5.2005
R2057 VSS.n338 VSS.n337 5.2005
R2058 VSS.n1596 VSS.n1595 5.2005
R2059 VSS.n1597 VSS.n1596 5.2005
R2060 VSS.n336 VSS.n335 5.2005
R2061 VSS.n1598 VSS.n336 5.2005
R2062 VSS.n1601 VSS.n1600 5.2005
R2063 VSS.n1600 VSS.n1599 5.2005
R2064 VSS.n1602 VSS.n334 5.2005
R2065 VSS.n334 VSS.n333 5.2005
R2066 VSS.n1604 VSS.n1603 5.2005
R2067 VSS.n1605 VSS.n1604 5.2005
R2068 VSS.n332 VSS.n331 5.2005
R2069 VSS.n1606 VSS.n332 5.2005
R2070 VSS.n1609 VSS.n1608 5.2005
R2071 VSS.n1608 VSS.n1607 5.2005
R2072 VSS.n1429 VSS.n330 5.2005
R2073 VSS.n1430 VSS.n1429 5.2005
R2074 VSS.n1428 VSS.n1427 5.2005
R2075 VSS.n1431 VSS.n1428 5.2005
R2076 VSS.n1434 VSS.n1433 5.2005
R2077 VSS.n1433 VSS.n1432 5.2005
R2078 VSS.n1435 VSS.n1426 5.2005
R2079 VSS.n1426 VSS.n1425 5.2005
R2080 VSS.n1437 VSS.n1436 5.2005
R2081 VSS.n1438 VSS.n1437 5.2005
R2082 VSS.n1424 VSS.n1423 5.2005
R2083 VSS.n1439 VSS.n1424 5.2005
R2084 VSS.n1442 VSS.n1441 5.2005
R2085 VSS.n1441 VSS.n1440 5.2005
R2086 VSS.n1443 VSS.n1422 5.2005
R2087 VSS.n1422 VSS.n1421 5.2005
R2088 VSS.n1445 VSS.n1444 5.2005
R2089 VSS.n1446 VSS.n1445 5.2005
R2090 VSS.n1420 VSS.n1419 5.2005
R2091 VSS.n1447 VSS.n1420 5.2005
R2092 VSS.n1451 VSS.n1450 5.2005
R2093 VSS.n1450 VSS.n1449 5.2005
R2094 VSS.n1452 VSS.n1418 5.2005
R2095 VSS.n1418 VSS.n1417 5.2005
R2096 VSS.n1454 VSS.n1453 5.2005
R2097 VSS.n1455 VSS.n1454 5.2005
R2098 VSS.n1416 VSS.n1415 5.2005
R2099 VSS.n1456 VSS.n1416 5.2005
R2100 VSS.n1459 VSS.n1458 5.2005
R2101 VSS.n1458 VSS.n1457 5.2005
R2102 VSS.n1460 VSS.n1414 5.2005
R2103 VSS.n1414 VSS.n1413 5.2005
R2104 VSS.n1462 VSS.n1461 5.2005
R2105 VSS.n1463 VSS.n1462 5.2005
R2106 VSS.n1412 VSS.n1411 5.2005
R2107 VSS.n1464 VSS.n1412 5.2005
R2108 VSS.n1467 VSS.n1466 5.2005
R2109 VSS.n1466 VSS.n1465 5.2005
R2110 VSS.n1410 VSS.n1409 5.2005
R2111 VSS.n1409 VSS.n470 5.2005
R2112 VSS.n1408 VSS.n485 5.2005
R2113 VSS.n1408 VSS.n1407 5.2005
R2114 VSS.n1401 VSS.n486 5.2005
R2115 VSS.n1406 VSS.n486 5.2005
R2116 VSS.n1403 VSS.n1402 5.2005
R2117 VSS.n1404 VSS.n1403 5.2005
R2118 VSS.n1400 VSS.n490 5.2005
R2119 VSS.n490 VSS.n489 5.2005
R2120 VSS.n1399 VSS.n1398 5.2005
R2121 VSS.n1398 VSS.n1397 5.2005
R2122 VSS.n492 VSS.n491 5.2005
R2123 VSS.n1396 VSS.n492 5.2005
R2124 VSS.n1394 VSS.n1393 5.2005
R2125 VSS.n1395 VSS.n1394 5.2005
R2126 VSS.n1392 VSS.n494 5.2005
R2127 VSS.n494 VSS.n493 5.2005
R2128 VSS.n1391 VSS.n1390 5.2005
R2129 VSS.n1390 VSS.n1389 5.2005
R2130 VSS.n496 VSS.n495 5.2005
R2131 VSS.n497 VSS.n496 5.2005
R2132 VSS.n1291 VSS.n1290 5.2005
R2133 VSS.n1290 VSS.n1289 5.2005
R2134 VSS.n1293 VSS.n1292 5.2005
R2135 VSS.n1294 VSS.n1293 5.2005
R2136 VSS.n1288 VSS.n1287 5.2005
R2137 VSS.n1295 VSS.n1288 5.2005
R2138 VSS.n1298 VSS.n1297 5.2005
R2139 VSS.n1297 VSS.n1296 5.2005
R2140 VSS.n1299 VSS.n1286 5.2005
R2141 VSS.n1286 VSS.n1285 5.2005
R2142 VSS.n1301 VSS.n1300 5.2005
R2143 VSS.n1302 VSS.n1301 5.2005
R2144 VSS.n1284 VSS.n1283 5.2005
R2145 VSS.n1303 VSS.n1284 5.2005
R2146 VSS.n1306 VSS.n1305 5.2005
R2147 VSS.n1305 VSS.n1304 5.2005
R2148 VSS.n1282 VSS.n1281 5.2005
R2149 VSS.n1281 VSS.n523 5.2005
R2150 VSS.n1280 VSS.n538 5.2005
R2151 VSS.n1280 VSS.n1279 5.2005
R2152 VSS.n1273 VSS.n539 5.2005
R2153 VSS.n1278 VSS.n539 5.2005
R2154 VSS.n1275 VSS.n1274 5.2005
R2155 VSS.n1276 VSS.n1275 5.2005
R2156 VSS.n1272 VSS.n543 5.2005
R2157 VSS.n543 VSS.n542 5.2005
R2158 VSS.n1271 VSS.n1270 5.2005
R2159 VSS.n1270 VSS.n1269 5.2005
R2160 VSS.n545 VSS.n544 5.2005
R2161 VSS.n1268 VSS.n545 5.2005
R2162 VSS.n1266 VSS.n1265 5.2005
R2163 VSS.n1267 VSS.n1266 5.2005
R2164 VSS.n1264 VSS.n547 5.2005
R2165 VSS.n547 VSS.n546 5.2005
R2166 VSS.n1263 VSS.n1262 5.2005
R2167 VSS.n1262 VSS.n1261 5.2005
R2168 VSS.n549 VSS.n548 5.2005
R2169 VSS.n550 VSS.n549 5.2005
R2170 VSS.n1163 VSS.n1162 5.2005
R2171 VSS.n1162 VSS.n1161 5.2005
R2172 VSS.n1165 VSS.n1164 5.2005
R2173 VSS.n1166 VSS.n1165 5.2005
R2174 VSS.n1160 VSS.n1159 5.2005
R2175 VSS.n1167 VSS.n1160 5.2005
R2176 VSS.n1170 VSS.n1169 5.2005
R2177 VSS.n1169 VSS.n1168 5.2005
R2178 VSS.n1171 VSS.n1158 5.2005
R2179 VSS.n1158 VSS.n1157 5.2005
R2180 VSS.n1173 VSS.n1172 5.2005
R2181 VSS.n1174 VSS.n1173 5.2005
R2182 VSS.n1156 VSS.n1155 5.2005
R2183 VSS.n1175 VSS.n1156 5.2005
R2184 VSS.n1178 VSS.n1177 5.2005
R2185 VSS.n1177 VSS.n1176 5.2005
R2186 VSS.n1154 VSS.n1153 5.2005
R2187 VSS.n1153 VSS.n577 5.2005
R2188 VSS.n1152 VSS.n592 5.2005
R2189 VSS.n1152 VSS.n1151 5.2005
R2190 VSS.n1145 VSS.n593 5.2005
R2191 VSS.n1150 VSS.n593 5.2005
R2192 VSS.n1147 VSS.n1146 5.2005
R2193 VSS.n1148 VSS.n1147 5.2005
R2194 VSS.n1144 VSS.n597 5.2005
R2195 VSS.n597 VSS.n596 5.2005
R2196 VSS.n1143 VSS.n1142 5.2005
R2197 VSS.n1142 VSS.n1141 5.2005
R2198 VSS.n599 VSS.n598 5.2005
R2199 VSS.n1140 VSS.n599 5.2005
R2200 VSS.n1138 VSS.n1137 5.2005
R2201 VSS.n1139 VSS.n1138 5.2005
R2202 VSS.n1136 VSS.n601 5.2005
R2203 VSS.n601 VSS.n600 5.2005
R2204 VSS.n1135 VSS.n1134 5.2005
R2205 VSS.n1134 VSS.n1133 5.2005
R2206 VSS.n603 VSS.n602 5.2005
R2207 VSS.n604 VSS.n603 5.2005
R2208 VSS.n1074 VSS.n1073 5.2005
R2209 VSS.n1075 VSS.n1074 5.2005
R2210 VSS.n1078 VSS.n1077 5.2005
R2211 VSS.n1077 VSS.n1076 5.2005
R2212 VSS.n1079 VSS.n1072 5.2005
R2213 VSS.n1072 VSS.n1071 5.2005
R2214 VSS.n1081 VSS.n1080 5.2005
R2215 VSS.n1082 VSS.n1081 5.2005
R2216 VSS.n1069 VSS.n1068 5.2005
R2217 VSS.n1083 VSS.n1069 5.2005
R2218 VSS.n1086 VSS.n1085 5.2005
R2219 VSS.n1085 VSS.n1084 5.2005
R2220 VSS.n1087 VSS.n622 5.2005
R2221 VSS.n1070 VSS.n622 5.2005
R2222 VSS.n1089 VSS.n1088 5.2005
R2223 VSS.n1090 VSS.n1089 5.2005
R2224 VSS.n2134 VSS.n168 5.2005
R2225 VSS.n2137 VSS.n2135 5.2005
R2226 VSS.n2140 VSS.n2139 5.2005
R2227 VSS.n2141 VSS.n2133 5.2005
R2228 VSS.n2143 VSS.n2142 5.2005
R2229 VSS.n2145 VSS.n2132 5.2005
R2230 VSS.n2148 VSS.n2147 5.2005
R2231 VSS.n2149 VSS.n2131 5.2005
R2232 VSS.n2151 VSS.n2150 5.2005
R2233 VSS.n2153 VSS.n2130 5.2005
R2234 VSS.n2156 VSS.n2155 5.2005
R2235 VSS.n2157 VSS.n2129 5.2005
R2236 VSS.n2159 VSS.n2158 5.2005
R2237 VSS.n2161 VSS.n2126 5.2005
R2238 VSS.n2164 VSS.n2163 5.2005
R2239 VSS.n2165 VSS.n2125 5.2005
R2240 VSS.n2167 VSS.n2166 5.2005
R2241 VSS.n2169 VSS.n2124 5.2005
R2242 VSS.n2171 VSS.n2170 5.2005
R2243 VSS.n2173 VSS.n2172 5.2005
R2244 VSS.n2174 VSS.n2122 5.2005
R2245 VSS.n2177 VSS.n2176 5.2005
R2246 VSS.n2183 VSS.n55 5.2005
R2247 VSS.n2183 VSS.n2182 5.2005
R2248 VSS.n2186 VSS.n2185 5.2005
R2249 VSS.n2187 VSS.n2186 5.2005
R2250 VSS.n2184 VSS.n167 5.2005
R2251 VSS.n167 VSS.n165 5.2005
R2252 VSS.n157 VSS.n156 5.2005
R2253 VSS.n159 VSS.n157 5.2005
R2254 VSS.n2197 VSS.n2196 5.2005
R2255 VSS.n2196 VSS.n2195 5.2005
R2256 VSS.n2198 VSS.n153 5.2005
R2257 VSS.n2127 VSS.n153 5.2005
R2258 VSS.n2200 VSS.n2199 5.2005
R2259 VSS.n2201 VSS.n2200 5.2005
R2260 VSS.n155 VSS.n152 5.2005
R2261 VSS.n152 VSS.n150 5.2005
R2262 VSS.n154 VSS.n143 5.2005
R2263 VSS.n2102 VSS.n143 5.2005
R2264 VSS.n2210 VSS.n144 5.2005
R2265 VSS.n2210 VSS.n2209 5.2005
R2266 VSS.n2211 VSS.n141 5.2005
R2267 VSS.n2214 VSS.n2213 5.2005
R2268 VSS.n2215 VSS.n138 5.2005
R2269 VSS.n2217 VSS.n2216 5.2005
R2270 VSS.n2218 VSS.n2217 5.2005
R2271 VSS.n140 VSS.n137 5.2005
R2272 VSS.n137 VSS.n135 5.2005
R2273 VSS.n139 VSS.n128 5.2005
R2274 VSS.n130 VSS.n128 5.2005
R2275 VSS.n2227 VSS.n129 5.2005
R2276 VSS.n2227 VSS.n2226 5.2005
R2277 VSS.n2228 VSS.n57 5.2005
R2278 VSS.n2229 VSS.n2228 5.2005
R2279 VSS.n60 VSS.n56 5.2005
R2280 VSS.n1926 VSS.n60 5.2005
R2281 VSS.n1921 VSS.n1920 5.2005
R2282 VSS.n1924 VSS.n1921 5.2005
R2283 VSS.n1936 VSS.n1935 5.2005
R2284 VSS.n1935 VSS.n1934 5.2005
R2285 VSS.n1937 VSS.n1917 5.2005
R2286 VSS.n1922 VSS.n1917 5.2005
R2287 VSS.n1939 VSS.n1938 5.2005
R2288 VSS.n1940 VSS.n1939 5.2005
R2289 VSS.n1919 VSS.n1916 5.2005
R2290 VSS.n1916 VSS.n1914 5.2005
R2291 VSS.n1918 VSS.n225 5.2005
R2292 VSS.n229 VSS.n225 5.2005
R2293 VSS.n1949 VSS.n226 5.2005
R2294 VSS.n1949 VSS.n1948 5.2005
R2295 VSS.n1950 VSS.n54 5.2005
R2296 VSS.n1951 VSS.n1950 5.2005
R2297 VSS.n1900 VSS.n224 5.2005
R2298 VSS.n1906 VSS.n224 5.2005
R2299 VSS.n1902 VSS.n1901 5.2005
R2300 VSS.n1899 VSS.n1887 5.2005
R2301 VSS.n1898 VSS.n1897 5.2005
R2302 VSS.n1896 VSS.n1895 5.2005
R2303 VSS.n1894 VSS.n1888 5.2005
R2304 VSS.n1892 VSS.n1891 5.2005
R2305 VSS.n1890 VSS.n52 5.2005
R2306 VSS.n2289 VSS.n53 5.2005
R2307 VSS.n2289 VSS.n2288 5.2005
R2308 VSS.n2286 VSS.n51 5.2005
R2309 VSS.n2285 VSS.n2284 5.2005
R2310 VSS.n2283 VSS.n2282 5.2005
R2311 VSS.n2281 VSS.n2244 5.2005
R2312 VSS.n2279 VSS.n2278 5.2005
R2313 VSS.n2277 VSS.n2245 5.2005
R2314 VSS.n2276 VSS.n2275 5.2005
R2315 VSS.n2273 VSS.n2246 5.2005
R2316 VSS.n2267 VSS.n2247 5.2005
R2317 VSS.n2269 VSS.n2268 5.2005
R2318 VSS.n2266 VSS.n2248 5.2005
R2319 VSS.n2265 VSS.n2264 5.2005
R2320 VSS.n2264 VSS.n2263 5.2005
R2321 VSS.n2250 VSS.n2249 5.2005
R2322 VSS.n2262 VSS.n2250 5.2005
R2323 VSS.n2260 VSS.n2259 5.2005
R2324 VSS.n2261 VSS.n2260 5.2005
R2325 VSS.n2258 VSS.n2252 5.2005
R2326 VSS.n2252 VSS.n2251 5.2005
R2327 VSS.n2257 VSS.n2256 5.2005
R2328 VSS.n2256 VSS.n2255 5.2005
R2329 VSS.n2253 VSS.n3 5.2005
R2330 VSS.n2254 VSS.n2253 5.2005
R2331 VSS.n2358 VSS.n5 5.2005
R2332 VSS.n9 VSS.n5 5.2005
R2333 VSS.n2358 VSS.n2357 5.2005
R2334 VSS.n2357 VSS.n2356 5.2005
R2335 VSS.n6 VSS.n2 5.2005
R2336 VSS.n8 VSS.n6 5.2005
R2337 VSS.n1570 VSS.n1569 5.2005
R2338 VSS.n1571 VSS.n1570 5.2005
R2339 VSS.n1568 VSS.n352 5.2005
R2340 VSS.n352 VSS.n351 5.2005
R2341 VSS.n1567 VSS.n1566 5.2005
R2342 VSS.n1566 VSS.n1565 5.2005
R2343 VSS.n354 VSS.n353 5.2005
R2344 VSS.n1564 VSS.n354 5.2005
R2345 VSS.n1562 VSS.n1561 5.2005
R2346 VSS.n1563 VSS.n1562 5.2005
R2347 VSS.n1560 VSS.n356 5.2005
R2348 VSS.n356 VSS.n355 5.2005
R2349 VSS.n1559 VSS.n1558 5.2005
R2350 VSS.n1558 VSS.n1557 5.2005
R2351 VSS.n358 VSS.n357 5.2005
R2352 VSS.n1556 VSS.n358 5.2005
R2353 VSS.n1554 VSS.n1553 5.2005
R2354 VSS.n1555 VSS.n1554 5.2005
R2355 VSS.n1552 VSS.n360 5.2005
R2356 VSS.n360 VSS.n359 5.2005
R2357 VSS.n1551 VSS.n1550 5.2005
R2358 VSS.n1550 VSS.n1549 5.2005
R2359 VSS.n362 VSS.n361 5.2005
R2360 VSS.n1548 VSS.n362 5.2005
R2361 VSS.n1546 VSS.n1545 5.2005
R2362 VSS.n1547 VSS.n1546 5.2005
R2363 VSS.n1544 VSS.n364 5.2005
R2364 VSS.n364 VSS.n363 5.2005
R2365 VSS.n1543 VSS.n1542 5.2005
R2366 VSS.n1542 VSS.n1541 5.2005
R2367 VSS.n366 VSS.n365 5.2005
R2368 VSS.n1540 VSS.n366 5.2005
R2369 VSS.n1538 VSS.n1537 5.2005
R2370 VSS.n1539 VSS.n1538 5.2005
R2371 VSS.n1537 VSS.n1536 5.2005
R2372 VSS.n1536 VSS.n1535 5.2005
R2373 VSS.n424 VSS.n369 5.2005
R2374 VSS.n1534 VSS.n424 5.2005
R2375 VSS.n1532 VSS.n1531 5.2005
R2376 VSS.n1533 VSS.n1532 5.2005
R2377 VSS.n1530 VSS.n426 5.2005
R2378 VSS.n1526 VSS.n426 5.2005
R2379 VSS.n1529 VSS.n1528 5.2005
R2380 VSS.n1528 VSS.n1527 5.2005
R2381 VSS.n428 VSS.n427 5.2005
R2382 VSS.n1525 VSS.n428 5.2005
R2383 VSS.n1523 VSS.n1522 5.2005
R2384 VSS.n1524 VSS.n1523 5.2005
R2385 VSS.n1521 VSS.n430 5.2005
R2386 VSS.n430 VSS.n429 5.2005
R2387 VSS.n1520 VSS.n1519 5.2005
R2388 VSS.n1519 VSS.n1518 5.2005
R2389 VSS.n432 VSS.n431 5.2005
R2390 VSS.n1517 VSS.n432 5.2005
R2391 VSS.n1515 VSS.n1514 5.2005
R2392 VSS.n1516 VSS.n1515 5.2005
R2393 VSS.n435 VSS.n434 5.2005
R2394 VSS.n434 VSS.n433 5.2005
R2395 VSS.n451 VSS.n450 5.2005
R2396 VSS.n452 VSS.n451 5.2005
R2397 VSS.n448 VSS.n447 5.2005
R2398 VSS.n453 VSS.n448 5.2005
R2399 VSS.n456 VSS.n455 5.2005
R2400 VSS.n455 VSS.n454 5.2005
R2401 VSS.n457 VSS.n446 5.2005
R2402 VSS.n449 VSS.n446 5.2005
R2403 VSS.n459 VSS.n458 5.2005
R2404 VSS.n459 VSS.n445 5.2005
R2405 VSS.n460 VSS.n439 5.2005
R2406 VSS.n461 VSS.n460 5.2005
R2407 VSS.n1511 VSS.n441 5.2005
R2408 VSS.n462 VSS.n441 5.2005
R2409 VSS.n1511 VSS.n1510 5.2005
R2410 VSS.n1510 VSS.n1509 5.2005
R2411 VSS.n442 VSS.n438 5.2005
R2412 VSS.n444 VSS.n442 5.2005
R2413 VSS.n1370 VSS.n1369 5.2005
R2414 VSS.n1369 VSS.n488 5.2005
R2415 VSS.n1371 VSS.n1368 5.2005
R2416 VSS.n1368 VSS.n487 5.2005
R2417 VSS.n1373 VSS.n1372 5.2005
R2418 VSS.n1374 VSS.n1373 5.2005
R2419 VSS.n1367 VSS.n1366 5.2005
R2420 VSS.n1375 VSS.n1367 5.2005
R2421 VSS.n1378 VSS.n1377 5.2005
R2422 VSS.n1377 VSS.n1376 5.2005
R2423 VSS.n1379 VSS.n1365 5.2005
R2424 VSS.n1365 VSS.n1364 5.2005
R2425 VSS.n1381 VSS.n1380 5.2005
R2426 VSS.n1382 VSS.n1381 5.2005
R2427 VSS.n501 VSS.n499 5.2005
R2428 VSS.n1383 VSS.n501 5.2005
R2429 VSS.n1386 VSS.n1385 5.2005
R2430 VSS.n1385 VSS.n1384 5.2005
R2431 VSS.n500 VSS.n498 5.2005
R2432 VSS.n1363 VSS.n500 5.2005
R2433 VSS.n1361 VSS.n1360 5.2005
R2434 VSS.n1362 VSS.n1361 5.2005
R2435 VSS.n1359 VSS.n503 5.2005
R2436 VSS.n503 VSS.n502 5.2005
R2437 VSS.n1358 VSS.n1357 5.2005
R2438 VSS.n1357 VSS.n1356 5.2005
R2439 VSS.n505 VSS.n504 5.2005
R2440 VSS.n1355 VSS.n505 5.2005
R2441 VSS.n1353 VSS.n1352 5.2005
R2442 VSS.n1354 VSS.n1353 5.2005
R2443 VSS.n1351 VSS.n507 5.2005
R2444 VSS.n507 VSS.n506 5.2005
R2445 VSS.n1350 VSS.n510 5.2005
R2446 VSS.n515 VSS.n510 5.2005
R2447 VSS.n1350 VSS.n1349 5.2005
R2448 VSS.n1349 VSS.n1348 5.2005
R2449 VSS.n512 VSS.n508 5.2005
R2450 VSS.n514 VSS.n512 5.2005
R2451 VSS.n1242 VSS.n1241 5.2005
R2452 VSS.n1241 VSS.n541 5.2005
R2453 VSS.n1243 VSS.n1240 5.2005
R2454 VSS.n1240 VSS.n540 5.2005
R2455 VSS.n1245 VSS.n1244 5.2005
R2456 VSS.n1246 VSS.n1245 5.2005
R2457 VSS.n1239 VSS.n1238 5.2005
R2458 VSS.n1247 VSS.n1239 5.2005
R2459 VSS.n1250 VSS.n1249 5.2005
R2460 VSS.n1249 VSS.n1248 5.2005
R2461 VSS.n1251 VSS.n1237 5.2005
R2462 VSS.n1237 VSS.n1236 5.2005
R2463 VSS.n1253 VSS.n1252 5.2005
R2464 VSS.n1254 VSS.n1253 5.2005
R2465 VSS.n555 VSS.n552 5.2005
R2466 VSS.n1255 VSS.n555 5.2005
R2467 VSS.n1258 VSS.n1257 5.2005
R2468 VSS.n1257 VSS.n1256 5.2005
R2469 VSS.n554 VSS.n551 5.2005
R2470 VSS.n1235 VSS.n554 5.2005
R2471 VSS.n1233 VSS.n1232 5.2005
R2472 VSS.n1234 VSS.n1233 5.2005
R2473 VSS.n1231 VSS.n557 5.2005
R2474 VSS.n557 VSS.n556 5.2005
R2475 VSS.n1230 VSS.n1229 5.2005
R2476 VSS.n1229 VSS.n1228 5.2005
R2477 VSS.n559 VSS.n558 5.2005
R2478 VSS.n1227 VSS.n559 5.2005
R2479 VSS.n1225 VSS.n1224 5.2005
R2480 VSS.n1226 VSS.n1225 5.2005
R2481 VSS.n1223 VSS.n561 5.2005
R2482 VSS.n561 VSS.n560 5.2005
R2483 VSS.n1222 VSS.n564 5.2005
R2484 VSS.n569 VSS.n564 5.2005
R2485 VSS.n1222 VSS.n1221 5.2005
R2486 VSS.n1221 VSS.n1220 5.2005
R2487 VSS.n566 VSS.n562 5.2005
R2488 VSS.n568 VSS.n566 5.2005
R2489 VSS.n1114 VSS.n1113 5.2005
R2490 VSS.n1113 VSS.n595 5.2005
R2491 VSS.n1115 VSS.n1112 5.2005
R2492 VSS.n1112 VSS.n594 5.2005
R2493 VSS.n1117 VSS.n1116 5.2005
R2494 VSS.n1118 VSS.n1117 5.2005
R2495 VSS.n1111 VSS.n1110 5.2005
R2496 VSS.n1119 VSS.n1111 5.2005
R2497 VSS.n1122 VSS.n1121 5.2005
R2498 VSS.n1121 VSS.n1120 5.2005
R2499 VSS.n1123 VSS.n1109 5.2005
R2500 VSS.n1109 VSS.n1108 5.2005
R2501 VSS.n1125 VSS.n1124 5.2005
R2502 VSS.n1126 VSS.n1125 5.2005
R2503 VSS.n609 VSS.n606 5.2005
R2504 VSS.n1127 VSS.n609 5.2005
R2505 VSS.n1130 VSS.n1129 5.2005
R2506 VSS.n1129 VSS.n1128 5.2005
R2507 VSS.n608 VSS.n605 5.2005
R2508 VSS.n1107 VSS.n608 5.2005
R2509 VSS.n1105 VSS.n1104 5.2005
R2510 VSS.n1106 VSS.n1105 5.2005
R2511 VSS.n1103 VSS.n611 5.2005
R2512 VSS.n611 VSS.n610 5.2005
R2513 VSS.n1102 VSS.n1101 5.2005
R2514 VSS.n1101 VSS.n1100 5.2005
R2515 VSS.n613 VSS.n612 5.2005
R2516 VSS.n1099 VSS.n613 5.2005
R2517 VSS.n1097 VSS.n1096 5.2005
R2518 VSS.n1098 VSS.n1097 5.2005
R2519 VSS.n1095 VSS.n615 5.2005
R2520 VSS.n615 VSS.n614 5.2005
R2521 VSS.n1094 VSS.n1093 5.2005
R2522 VSS.n1093 VSS.n1092 5.2005
R2523 VSS.n96 VSS.n73 5.2005
R2524 VSS.n99 VSS.n98 5.2005
R2525 VSS.n100 VSS.n72 5.2005
R2526 VSS.n102 VSS.n101 5.2005
R2527 VSS.n104 VSS.n71 5.2005
R2528 VSS.n107 VSS.n106 5.2005
R2529 VSS.n108 VSS.n70 5.2005
R2530 VSS.n110 VSS.n109 5.2005
R2531 VSS.n112 VSS.n69 5.2005
R2532 VSS.n115 VSS.n114 5.2005
R2533 VSS.n116 VSS.n68 5.2005
R2534 VSS.n118 VSS.n117 5.2005
R2535 VSS.n120 VSS.n67 5.2005
R2536 VSS.n122 VSS.n121 5.2005
R2537 VSS.n121 VSS.n63 5.2005
R2538 VSS.n94 VSS.n93 5.2005
R2539 VSS.n80 VSS.n58 5.2005
R2540 VSS.n80 VSS.n63 5.2005
R2541 VSS.n83 VSS.n82 5.2005
R2542 VSS.n84 VSS.n79 5.2005
R2543 VSS.n86 VSS.n85 5.2005
R2544 VSS.n88 VSS.n78 5.2005
R2545 VSS.n91 VSS.n90 5.2005
R2546 VSS.n92 VSS.n74 5.2005
R2547 VSS.n2239 VSS.n59 5.2005
R2548 VSS.n126 VSS.n59 5.2005
R2549 VSS.n2239 VSS.n2238 5.2005
R2550 VSS.n2238 VSS.n2237 5.2005
R2551 VSS.n77 VSS.n75 4.55948
R2552 VSS.n2080 VSS.n180 4.5191
R2553 VSS.n77 VSS.n76 4.38259
R2554 VSS.n2164 VSS.n2128 3.87024
R2555 VSS.n2149 VSS.n2128 3.87024
R2556 VSS.n2120 VSS.n170 3.59261
R2557 VSS.n1997 VSS.n65 3.59261
R2558 VSS.n30 VSS.n28 3.59261
R2559 VSS.n1612 VSS.n328 3.59261
R2560 VSS.n483 VSS.n481 3.59261
R2561 VSS.n536 VSS.n534 3.59261
R2562 VSS.n590 VSS.n588 3.59261
R2563 VSS.n1065 VSS.n621 3.59261
R2564 VSS.n1792 VSS.n248 3.59261
R2565 VSS.t22 VSS.n206 3.52692
R2566 VSS.n2089 VSS.n2088 3.32459
R2567 VSS.n2092 VSS.n2091 3.32459
R2568 VSS.n2096 VSS.n177 3.32459
R2569 VSS.n2099 VSS.n2098 3.32459
R2570 VSS.n2108 VSS.n2107 3.32459
R2571 VSS.n2111 VSS.n2110 3.32459
R2572 VSS.n2116 VSS.n2115 3.32459
R2573 VSS.n2119 VSS.n2118 3.32459
R2574 VSS.n2010 VSS.n2009 3.32459
R2575 VSS.n2005 VSS.n1996 3.32459
R2576 VSS.n2003 VSS.n2002 3.32459
R2577 VSS.n1998 VSS.n1997 3.32459
R2578 VSS.n1698 VSS.n18 3.32459
R2579 VSS.n30 VSS.n19 3.32459
R2580 VSS.n1615 VSS.n326 3.32459
R2581 VSS.n1613 VSS.n1612 3.32459
R2582 VSS.n846 VSS.n471 3.32459
R2583 VSS.n483 VSS.n472 3.32459
R2584 VSS.n783 VSS.n524 3.32459
R2585 VSS.n536 VSS.n525 3.32459
R2586 VSS.n1022 VSS.n701 3.32459
R2587 VSS.n1018 VSS.n700 3.32459
R2588 VSS.n1014 VSS.n699 3.32459
R2589 VSS.n1010 VSS.n698 3.32459
R2590 VSS.n1006 VSS.n697 3.32459
R2591 VSS.n1002 VSS.n696 3.32459
R2592 VSS.n998 VSS.n578 3.32459
R2593 VSS.n590 VSS.n579 3.32459
R2594 VSS.n1005 VSS.n696 3.32459
R2595 VSS.n1009 VSS.n697 3.32459
R2596 VSS.n1013 VSS.n698 3.32459
R2597 VSS.n1017 VSS.n699 3.32459
R2598 VSS.n1021 VSS.n700 3.32459
R2599 VSS.n995 VSS.n701 3.32459
R2600 VSS.n673 VSS.n672 3.32459
R2601 VSS.n670 VSS.n624 3.32459
R2602 VSS.n666 VSS.n665 3.32459
R2603 VSS.n659 VSS.n626 3.32459
R2604 VSS.n658 VSS.n657 3.32459
R2605 VSS.n651 VSS.n628 3.32459
R2606 VSS.n650 VSS.n649 3.32459
R2607 VSS.n643 VSS.n630 3.32459
R2608 VSS.n641 VSS.n632 3.32459
R2609 VSS.n637 VSS.n636 3.32459
R2610 VSS.n589 VSS.n580 3.32459
R2611 VSS.n1201 VSS.n581 3.32459
R2612 VSS.n1197 VSS.n582 3.32459
R2613 VSS.n1193 VSS.n583 3.32459
R2614 VSS.n1189 VSS.n584 3.32459
R2615 VSS.n1185 VSS.n585 3.32459
R2616 VSS.n1181 VSS.n586 3.32459
R2617 VSS.n1209 VSS.n1208 3.32459
R2618 VSS.n1214 VSS.n572 3.32459
R2619 VSS.n571 VSS.n570 3.32459
R2620 VSS.n535 VSS.n526 3.32459
R2621 VSS.n1329 VSS.n527 3.32459
R2622 VSS.n1325 VSS.n528 3.32459
R2623 VSS.n1321 VSS.n529 3.32459
R2624 VSS.n1317 VSS.n530 3.32459
R2625 VSS.n1313 VSS.n531 3.32459
R2626 VSS.n1309 VSS.n532 3.32459
R2627 VSS.n1337 VSS.n1336 3.32459
R2628 VSS.n1342 VSS.n518 3.32459
R2629 VSS.n517 VSS.n516 3.32459
R2630 VSS.n482 VSS.n473 3.32459
R2631 VSS.n1490 VSS.n474 3.32459
R2632 VSS.n1486 VSS.n475 3.32459
R2633 VSS.n1482 VSS.n476 3.32459
R2634 VSS.n1478 VSS.n477 3.32459
R2635 VSS.n1474 VSS.n478 3.32459
R2636 VSS.n1470 VSS.n479 3.32459
R2637 VSS.n1498 VSS.n1497 3.32459
R2638 VSS.n1503 VSS.n465 3.32459
R2639 VSS.n464 VSS.n463 3.32459
R2640 VSS.n383 VSS.n382 3.32459
R2641 VSS.n388 VSS.n387 3.32459
R2642 VSS.n391 VSS.n390 3.32459
R2643 VSS.n396 VSS.n395 3.32459
R2644 VSS.n399 VSS.n398 3.32459
R2645 VSS.n404 VSS.n403 3.32459
R2646 VSS.n407 VSS.n406 3.32459
R2647 VSS.n412 VSS.n411 3.32459
R2648 VSS.n418 VSS.n371 3.32459
R2649 VSS.n421 VSS.n420 3.32459
R2650 VSS.n29 VSS.n20 3.32459
R2651 VSS.n2337 VSS.n21 3.32459
R2652 VSS.n2333 VSS.n22 3.32459
R2653 VSS.n2329 VSS.n23 3.32459
R2654 VSS.n2325 VSS.n24 3.32459
R2655 VSS.n2321 VSS.n25 3.32459
R2656 VSS.n2317 VSS.n26 3.32459
R2657 VSS.n2345 VSS.n2344 3.32459
R2658 VSS.n2350 VSS.n12 3.32459
R2659 VSS.n11 VSS.n10 3.32459
R2660 VSS.n2349 VSS.n11 3.32459
R2661 VSS.n14 VSS.n12 3.32459
R2662 VSS.n420 VSS.n419 3.32459
R2663 VSS.n415 VSS.n371 3.32459
R2664 VSS.n1502 VSS.n464 3.32459
R2665 VSS.n467 VSS.n465 3.32459
R2666 VSS.n1341 VSS.n517 3.32459
R2667 VSS.n520 VSS.n518 3.32459
R2668 VSS.n1213 VSS.n571 3.32459
R2669 VSS.n574 VSS.n572 3.32459
R2670 VSS.n638 VSS.n632 3.32459
R2671 VSS.n636 VSS.n635 3.32459
R2672 VSS.n997 VSS.n579 3.32459
R2673 VSS.n1001 VSS.n578 3.32459
R2674 VSS.n782 VSS.n525 3.32459
R2675 VSS.n786 VSS.n524 3.32459
R2676 VSS.n845 VSS.n472 3.32459
R2677 VSS.n849 VSS.n471 3.32459
R2678 VSS.n1614 VSS.n1613 3.32459
R2679 VSS.n326 VSS.n324 3.32459
R2680 VSS.n1697 VSS.n19 3.32459
R2681 VSS.n1701 VSS.n18 3.32459
R2682 VSS.n672 VSS.n671 3.32459
R2683 VSS.n667 VSS.n624 3.32459
R2684 VSS.n665 VSS.n664 3.32459
R2685 VSS.n660 VSS.n659 3.32459
R2686 VSS.n657 VSS.n656 3.32459
R2687 VSS.n652 VSS.n651 3.32459
R2688 VSS.n649 VSS.n648 3.32459
R2689 VSS.n644 VSS.n643 3.32459
R2690 VSS.n1208 VSS.n573 3.32459
R2691 VSS.n586 VSS.n576 3.32459
R2692 VSS.n1182 VSS.n585 3.32459
R2693 VSS.n1186 VSS.n584 3.32459
R2694 VSS.n1190 VSS.n583 3.32459
R2695 VSS.n1194 VSS.n582 3.32459
R2696 VSS.n1198 VSS.n581 3.32459
R2697 VSS.n1202 VSS.n580 3.32459
R2698 VSS.n1336 VSS.n519 3.32459
R2699 VSS.n532 VSS.n522 3.32459
R2700 VSS.n1310 VSS.n531 3.32459
R2701 VSS.n1314 VSS.n530 3.32459
R2702 VSS.n1318 VSS.n529 3.32459
R2703 VSS.n1322 VSS.n528 3.32459
R2704 VSS.n1326 VSS.n527 3.32459
R2705 VSS.n1330 VSS.n526 3.32459
R2706 VSS.n1497 VSS.n466 3.32459
R2707 VSS.n479 VSS.n469 3.32459
R2708 VSS.n1471 VSS.n478 3.32459
R2709 VSS.n1475 VSS.n477 3.32459
R2710 VSS.n1479 VSS.n476 3.32459
R2711 VSS.n1483 VSS.n475 3.32459
R2712 VSS.n1487 VSS.n474 3.32459
R2713 VSS.n1491 VSS.n473 3.32459
R2714 VSS.n413 VSS.n412 3.32459
R2715 VSS.n406 VSS.n374 3.32459
R2716 VSS.n405 VSS.n404 3.32459
R2717 VSS.n398 VSS.n376 3.32459
R2718 VSS.n397 VSS.n396 3.32459
R2719 VSS.n390 VSS.n378 3.32459
R2720 VSS.n389 VSS.n388 3.32459
R2721 VSS.n382 VSS.n380 3.32459
R2722 VSS.n2344 VSS.n13 3.32459
R2723 VSS.n26 VSS.n16 3.32459
R2724 VSS.n2318 VSS.n25 3.32459
R2725 VSS.n2322 VSS.n24 3.32459
R2726 VSS.n2326 VSS.n23 3.32459
R2727 VSS.n2330 VSS.n22 3.32459
R2728 VSS.n2334 VSS.n21 3.32459
R2729 VSS.n2338 VSS.n20 3.32459
R2730 VSS.n1999 VSS.n1998 3.32459
R2731 VSS.n2004 VSS.n2003 3.32459
R2732 VSS.n1996 VSS.n1994 3.32459
R2733 VSS.n2011 VSS.n2010 3.32459
R2734 VSS.n2093 VSS.n177 3.32459
R2735 VSS.n2091 VSS.n179 3.32459
R2736 VSS.n2089 VSS.n181 3.32459
R2737 VSS.n2098 VSS.n2097 3.32459
R2738 VSS.n2120 VSS.n2119 3.32459
R2739 VSS.n2117 VSS.n2116 3.32459
R2740 VSS.n2110 VSS.n173 3.32459
R2741 VSS.n2109 VSS.n2108 3.32459
R2742 VSS.n1061 VSS.n1060 3.32459
R2743 VSS.n1065 VSS.n1064 3.32459
R2744 VSS.n1062 VSS.n1061 3.32459
R2745 VSS.n1064 VSS.n1063 3.32459
R2746 VSS.n763 VSS.n762 3.32459
R2747 VSS.n760 VSS.n759 3.32459
R2748 VSS.n755 VSS.n744 3.32459
R2749 VSS.n753 VSS.n752 3.32459
R2750 VSS.n975 VSS.n974 3.32459
R2751 VSS.n970 VSS.n715 3.32459
R2752 VSS.n968 VSS.n967 3.32459
R2753 VSS.n963 VSS.n719 3.32459
R2754 VSS.n961 VSS.n960 3.32459
R2755 VSS.n955 VSS.n954 3.32459
R2756 VSS.n950 VSS.n817 3.32459
R2757 VSS.n948 VSS.n947 3.32459
R2758 VSS.n943 VSS.n820 3.32459
R2759 VSS.n940 VSS.n939 3.32459
R2760 VSS.n935 VSS.n825 3.32459
R2761 VSS.n933 VSS.n932 3.32459
R2762 VSS.n928 VSS.n829 3.32459
R2763 VSS.n926 VSS.n925 3.32459
R2764 VSS.n920 VSS.n919 3.32459
R2765 VSS.n915 VSS.n880 3.32459
R2766 VSS.n913 VSS.n912 3.32459
R2767 VSS.n908 VSS.n883 3.32459
R2768 VSS.n905 VSS.n904 3.32459
R2769 VSS.n900 VSS.n291 3.32459
R2770 VSS.n896 VSS.n292 3.32459
R2771 VSS.n892 VSS.n293 3.32459
R2772 VSS.n887 VSS.n294 3.32459
R2773 VSS.n299 VSS.n295 3.32459
R2774 VSS.n297 VSS.n296 3.32459
R2775 VSS.n305 VSS.n290 3.32459
R2776 VSS.n1647 VSS.n288 3.32459
R2777 VSS.n1656 VSS.n1655 3.32459
R2778 VSS.n1660 VSS.n275 3.32459
R2779 VSS.n1664 VSS.n276 3.32459
R2780 VSS.n1668 VSS.n277 3.32459
R2781 VSS.n1672 VSS.n278 3.32459
R2782 VSS.n1680 VSS.n279 3.32459
R2783 VSS.n1676 VSS.n280 3.32459
R2784 VSS.n281 VSS.n274 3.32459
R2785 VSS.n1730 VSS.n272 3.32459
R2786 VSS.n1739 VSS.n1738 3.32459
R2787 VSS.n1740 VSS.n269 3.32459
R2788 VSS.n1747 VSS.n1746 3.32459
R2789 VSS.n1748 VSS.n267 3.32459
R2790 VSS.n1755 VSS.n1754 3.32459
R2791 VSS.n1979 VSS.n1978 3.32459
R2792 VSS.n1976 VSS.n1975 3.32459
R2793 VSS.n1971 VSS.n222 3.32459
R2794 VSS.n1969 VSS.n1968 3.32459
R2795 VSS.n1964 VSS.n1956 3.32459
R2796 VSS.n1962 VSS.n1961 3.32459
R2797 VSS.n1957 VSS.n213 3.32459
R2798 VSS.n2055 VSS.n212 3.32459
R2799 VSS.n2050 VSS.n211 3.32459
R2800 VSS.n2044 VSS.n210 3.32459
R2801 VSS.n2040 VSS.n209 3.32459
R2802 VSS.n2036 VSS.n208 3.32459
R2803 VSS.n2033 VSS.n195 3.32459
R2804 VSS.n2034 VSS.n2033 3.32459
R2805 VSS.n2039 VSS.n208 3.32459
R2806 VSS.n2043 VSS.n209 3.32459
R2807 VSS.n2048 VSS.n210 3.32459
R2808 VSS.n2054 VSS.n211 3.32459
R2809 VSS.n214 VSS.n212 3.32459
R2810 VSS.n1958 VSS.n1957 3.32459
R2811 VSS.n1963 VSS.n1962 3.32459
R2812 VSS.n1956 VSS.n1954 3.32459
R2813 VSS.n1970 VSS.n1969 3.32459
R2814 VSS.n222 VSS.n220 3.32459
R2815 VSS.n1977 VSS.n1976 3.32459
R2816 VSS.n1980 VSS.n1979 3.32459
R2817 VSS.n1754 VSS.n1753 3.32459
R2818 VSS.n1749 VSS.n1748 3.32459
R2819 VSS.n1746 VSS.n1745 3.32459
R2820 VSS.n1741 VSS.n1740 3.32459
R2821 VSS.n1738 VSS.n271 3.32459
R2822 VSS.n1731 VSS.n1730 3.32459
R2823 VSS.n1675 VSS.n281 3.32459
R2824 VSS.n1679 VSS.n280 3.32459
R2825 VSS.n1683 VSS.n279 3.32459
R2826 VSS.n1669 VSS.n278 3.32459
R2827 VSS.n1665 VSS.n277 3.32459
R2828 VSS.n1661 VSS.n276 3.32459
R2829 VSS.n1657 VSS.n275 3.32459
R2830 VSS.n1655 VSS.n287 3.32459
R2831 VSS.n1648 VSS.n1647 3.32459
R2832 VSS.n305 VSS.n304 3.32459
R2833 VSS.n300 VSS.n296 3.32459
R2834 VSS.n309 VSS.n295 3.32459
R2835 VSS.n891 VSS.n294 3.32459
R2836 VSS.n895 VSS.n293 3.32459
R2837 VSS.n899 VSS.n292 3.32459
R2838 VSS.n885 VSS.n291 3.32459
R2839 VSS.n905 VSS.n884 3.32459
R2840 VSS.n883 VSS.n881 3.32459
R2841 VSS.n914 VSS.n913 3.32459
R2842 VSS.n880 VSS.n878 3.32459
R2843 VSS.n921 VSS.n920 3.32459
R2844 VSS.n927 VSS.n926 3.32459
R2845 VSS.n829 VSS.n827 3.32459
R2846 VSS.n934 VSS.n933 3.32459
R2847 VSS.n825 VSS.n822 3.32459
R2848 VSS.n940 VSS.n821 3.32459
R2849 VSS.n820 VSS.n818 3.32459
R2850 VSS.n949 VSS.n948 3.32459
R2851 VSS.n817 VSS.n815 3.32459
R2852 VSS.n956 VSS.n955 3.32459
R2853 VSS.n962 VSS.n961 3.32459
R2854 VSS.n719 VSS.n717 3.32459
R2855 VSS.n969 VSS.n968 3.32459
R2856 VSS.n715 VSS.n713 3.32459
R2857 VSS.n975 VSS.n712 3.32459
R2858 VSS.n754 VSS.n753 3.32459
R2859 VSS.n744 VSS.n742 3.32459
R2860 VSS.n761 VSS.n760 3.32459
R2861 VSS.n764 VSS.n763 3.32459
R2862 VSS.n1800 VSS.n1797 3.32459
R2863 VSS.n1807 VSS.n1806 3.32459
R2864 VSS.n1811 VSS.n1795 3.32459
R2865 VSS.n1814 VSS.n1813 3.32459
R2866 VSS.n1831 VSS.n1830 3.32459
R2867 VSS.n1828 VSS.n1827 3.32459
R2868 VSS.n1823 VSS.n1820 3.32459
R2869 VSS.n200 VSS.n145 3.32459
R2870 VSS.n201 VSS.n200 3.32459
R2871 VSS.n1820 VSS.n1818 3.32459
R2872 VSS.n1829 VSS.n1828 3.32459
R2873 VSS.n1832 VSS.n1831 3.32459
R2874 VSS.n1813 VSS.n1812 3.32459
R2875 VSS.n1808 VSS.n1795 3.32459
R2876 VSS.n1806 VSS.n1805 3.32459
R2877 VSS.n1801 VSS.n1800 3.32459
R2878 VSS.n2176 VSS.n2175 3.32459
R2879 VSS.n2173 VSS.n2123 3.32459
R2880 VSS.n2169 VSS.n2168 3.32459
R2881 VSS.n2162 VSS.n2125 3.32459
R2882 VSS.n2161 VSS.n2160 3.32459
R2883 VSS.n2154 VSS.n2129 3.32459
R2884 VSS.n2153 VSS.n2152 3.32459
R2885 VSS.n2146 VSS.n2131 3.32459
R2886 VSS.n2145 VSS.n2144 3.32459
R2887 VSS.n2138 VSS.n2133 3.32459
R2888 VSS.n2137 VSS.n2136 3.32459
R2889 VSS.n2136 VSS.n168 3.32459
R2890 VSS.n2139 VSS.n2138 3.32459
R2891 VSS.n2144 VSS.n2143 3.32459
R2892 VSS.n2147 VSS.n2146 3.32459
R2893 VSS.n2152 VSS.n2151 3.32459
R2894 VSS.n2155 VSS.n2154 3.32459
R2895 VSS.n2160 VSS.n2159 3.32459
R2896 VSS.n2163 VSS.n2162 3.32459
R2897 VSS.n2168 VSS.n2167 3.32459
R2898 VSS.n2170 VSS.n2123 3.32459
R2899 VSS.n2175 VSS.n2174 3.32459
R2900 VSS.n2270 VSS.n2269 3.32459
R2901 VSS.n2273 VSS.n2272 3.32459
R2902 VSS.n2274 VSS.n2245 3.32459
R2903 VSS.n2281 VSS.n2280 3.32459
R2904 VSS.n2285 VSS.n2243 3.32459
R2905 VSS.n2288 VSS.n2287 3.32459
R2906 VSS.n1890 VSS.n1889 3.32459
R2907 VSS.n1894 VSS.n1893 3.32459
R2908 VSS.n1897 VSS.n235 3.32459
R2909 VSS.n2212 VSS.n2211 3.32459
R2910 VSS.n2213 VSS.n2212 3.32459
R2911 VSS.n1895 VSS.n235 3.32459
R2912 VSS.n1893 VSS.n1892 3.32459
R2913 VSS.n1889 VSS.n53 3.32459
R2914 VSS.n2287 VSS.n2286 3.32459
R2915 VSS.n2282 VSS.n2243 3.32459
R2916 VSS.n2280 VSS.n2279 3.32459
R2917 VSS.n2275 VSS.n2274 3.32459
R2918 VSS.n2272 VSS.n2247 3.32459
R2919 VSS.n2270 VSS.n2248 3.32459
R2920 VSS.n120 VSS.n119 3.32459
R2921 VSS.n113 VSS.n68 3.32459
R2922 VSS.n112 VSS.n111 3.32459
R2923 VSS.n105 VSS.n70 3.32459
R2924 VSS.n104 VSS.n103 3.32459
R2925 VSS.n97 VSS.n72 3.32459
R2926 VSS.n96 VSS.n95 3.32459
R2927 VSS.n89 VSS.n74 3.32459
R2928 VSS.n88 VSS.n87 3.32459
R2929 VSS.n81 VSS.n79 3.32459
R2930 VSS.n98 VSS.n97 3.32459
R2931 VSS.n103 VSS.n102 3.32459
R2932 VSS.n106 VSS.n105 3.32459
R2933 VSS.n111 VSS.n110 3.32459
R2934 VSS.n114 VSS.n113 3.32459
R2935 VSS.n119 VSS.n118 3.32459
R2936 VSS.n95 VSS.n94 3.32459
R2937 VSS.n82 VSS.n81 3.32459
R2938 VSS.n87 VSS.n86 3.32459
R2939 VSS.n90 VSS.n89 3.32459
R2940 VSS.n93 VSS.n77 1.95679
R2941 VSS.n2240 VSS.n55 1.4552
R2942 VSS.n766 VSS 1.33138
R2943 VSS.n2046 VSS.n184 1.32688
R2944 VSS.n2052 VSS.n1982 1.316
R2945 VSS.n1682 VSS.n266 1.316
R2946 VSS.n1671 VSS.n285 1.316
R2947 VSS.n889 VSS.n877 1.316
R2948 VSS.n831 VSS.n814 1.316
R2949 VSS.n767 VSS.n766 1.316
R2950 VSS.n1027 VSS.n696 0.939203
R2951 VSS.n1027 VSS.n697 0.939203
R2952 VSS.n1027 VSS.n698 0.939203
R2953 VSS.n1027 VSS.n699 0.939203
R2954 VSS.n1027 VSS.n700 0.939203
R2955 VSS.n1027 VSS.n701 0.939203
R2956 VSS.n2355 VSS.n11 0.939203
R2957 VSS.n2355 VSS.n12 0.939203
R2958 VSS.n420 VSS.n367 0.939203
R2959 VSS.n371 VSS.n367 0.939203
R2960 VSS.n1508 VSS.n464 0.939203
R2961 VSS.n1508 VSS.n465 0.939203
R2962 VSS.n1347 VSS.n517 0.939203
R2963 VSS.n1347 VSS.n518 0.939203
R2964 VSS.n1219 VSS.n571 0.939203
R2965 VSS.n1219 VSS.n572 0.939203
R2966 VSS.n632 VSS.n618 0.939203
R2967 VSS.n636 VSS.n618 0.939203
R2968 VSS.n1207 VSS.n579 0.939203
R2969 VSS.n1207 VSS.n578 0.939203
R2970 VSS.n1335 VSS.n525 0.939203
R2971 VSS.n1335 VSS.n524 0.939203
R2972 VSS.n1496 VSS.n472 0.939203
R2973 VSS.n1496 VSS.n471 0.939203
R2974 VSS.n1613 VSS.n327 0.939203
R2975 VSS.n327 VSS.n326 0.939203
R2976 VSS.n2343 VSS.n19 0.939203
R2977 VSS.n2343 VSS.n18 0.939203
R2978 VSS.n672 VSS.n619 0.939203
R2979 VSS.n624 VSS.n619 0.939203
R2980 VSS.n665 VSS.n619 0.939203
R2981 VSS.n659 VSS.n619 0.939203
R2982 VSS.n657 VSS.n619 0.939203
R2983 VSS.n651 VSS.n619 0.939203
R2984 VSS.n649 VSS.n619 0.939203
R2985 VSS.n643 VSS.n619 0.939203
R2986 VSS.n1208 VSS.n1207 0.939203
R2987 VSS.n1207 VSS.n586 0.939203
R2988 VSS.n1207 VSS.n585 0.939203
R2989 VSS.n1207 VSS.n584 0.939203
R2990 VSS.n1207 VSS.n583 0.939203
R2991 VSS.n1207 VSS.n582 0.939203
R2992 VSS.n1207 VSS.n581 0.939203
R2993 VSS.n1207 VSS.n580 0.939203
R2994 VSS.n1336 VSS.n1335 0.939203
R2995 VSS.n1335 VSS.n532 0.939203
R2996 VSS.n1335 VSS.n531 0.939203
R2997 VSS.n1335 VSS.n530 0.939203
R2998 VSS.n1335 VSS.n529 0.939203
R2999 VSS.n1335 VSS.n528 0.939203
R3000 VSS.n1335 VSS.n527 0.939203
R3001 VSS.n1335 VSS.n526 0.939203
R3002 VSS.n1497 VSS.n1496 0.939203
R3003 VSS.n1496 VSS.n479 0.939203
R3004 VSS.n1496 VSS.n478 0.939203
R3005 VSS.n1496 VSS.n477 0.939203
R3006 VSS.n1496 VSS.n476 0.939203
R3007 VSS.n1496 VSS.n475 0.939203
R3008 VSS.n1496 VSS.n474 0.939203
R3009 VSS.n1496 VSS.n473 0.939203
R3010 VSS.n412 VSS.n327 0.939203
R3011 VSS.n406 VSS.n327 0.939203
R3012 VSS.n404 VSS.n327 0.939203
R3013 VSS.n398 VSS.n327 0.939203
R3014 VSS.n396 VSS.n327 0.939203
R3015 VSS.n390 VSS.n327 0.939203
R3016 VSS.n388 VSS.n327 0.939203
R3017 VSS.n382 VSS.n327 0.939203
R3018 VSS.n2344 VSS.n2343 0.939203
R3019 VSS.n2343 VSS.n26 0.939203
R3020 VSS.n2343 VSS.n25 0.939203
R3021 VSS.n2343 VSS.n24 0.939203
R3022 VSS.n2343 VSS.n23 0.939203
R3023 VSS.n2343 VSS.n22 0.939203
R3024 VSS.n2343 VSS.n21 0.939203
R3025 VSS.n2343 VSS.n20 0.939203
R3026 VSS.n1998 VSS.n63 0.939203
R3027 VSS.n2003 VSS.n63 0.939203
R3028 VSS.n1996 VSS.n63 0.939203
R3029 VSS.n2010 VSS.n63 0.939203
R3030 VSS.n2090 VSS.n177 0.939203
R3031 VSS.n2091 VSS.n2090 0.939203
R3032 VSS.n2090 VSS.n2089 0.939203
R3033 VSS.n2098 VSS.n169 0.939203
R3034 VSS.n2119 VSS.n169 0.939203
R3035 VSS.n2116 VSS.n169 0.939203
R3036 VSS.n2110 VSS.n169 0.939203
R3037 VSS.n2108 VSS.n169 0.939203
R3038 VSS.n1061 VSS.n619 0.939203
R3039 VSS.n1064 VSS.n619 0.939203
R3040 VSS.n2033 VSS.n196 0.939203
R3041 VSS.n2060 VSS.n208 0.939203
R3042 VSS.n2060 VSS.n209 0.939203
R3043 VSS.n2060 VSS.n210 0.939203
R3044 VSS.n2060 VSS.n211 0.939203
R3045 VSS.n2060 VSS.n212 0.939203
R3046 VSS.n1957 VSS.n199 0.939203
R3047 VSS.n1962 VSS.n199 0.939203
R3048 VSS.n1956 VSS.n1953 0.939203
R3049 VSS.n1969 VSS.n1953 0.939203
R3050 VSS.n1953 VSS.n222 0.939203
R3051 VSS.n1976 VSS.n218 0.939203
R3052 VSS.n1979 VSS.n218 0.939203
R3053 VSS.n1754 VSS.n218 0.939203
R3054 VSS.n1748 VSS.n218 0.939203
R3055 VSS.n1746 VSS.n218 0.939203
R3056 VSS.n1740 VSS.n218 0.939203
R3057 VSS.n1738 VSS.n1737 0.939203
R3058 VSS.n1730 VSS.n1729 0.939203
R3059 VSS.n1729 VSS.n281 0.939203
R3060 VSS.n1729 VSS.n280 0.939203
R3061 VSS.n1729 VSS.n279 0.939203
R3062 VSS.n1729 VSS.n278 0.939203
R3063 VSS.n1729 VSS.n277 0.939203
R3064 VSS.n1729 VSS.n276 0.939203
R3065 VSS.n1729 VSS.n275 0.939203
R3066 VSS.n1655 VSS.n1654 0.939203
R3067 VSS.n1647 VSS.n1646 0.939203
R3068 VSS.n1646 VSS.n305 0.939203
R3069 VSS.n1646 VSS.n296 0.939203
R3070 VSS.n1646 VSS.n295 0.939203
R3071 VSS.n1646 VSS.n294 0.939203
R3072 VSS.n1646 VSS.n293 0.939203
R3073 VSS.n1646 VSS.n292 0.939203
R3074 VSS.n1646 VSS.n291 0.939203
R3075 VSS.n906 VSS.n905 0.939203
R3076 VSS.n883 VSS.n826 0.939203
R3077 VSS.n913 VSS.n826 0.939203
R3078 VSS.n880 VSS.n826 0.939203
R3079 VSS.n920 VSS.n826 0.939203
R3080 VSS.n926 VSS.n826 0.939203
R3081 VSS.n829 VSS.n826 0.939203
R3082 VSS.n933 VSS.n826 0.939203
R3083 VSS.n826 VSS.n825 0.939203
R3084 VSS.n941 VSS.n940 0.939203
R3085 VSS.n820 VSS.n716 0.939203
R3086 VSS.n948 VSS.n716 0.939203
R3087 VSS.n817 VSS.n716 0.939203
R3088 VSS.n955 VSS.n716 0.939203
R3089 VSS.n961 VSS.n716 0.939203
R3090 VSS.n719 VSS.n716 0.939203
R3091 VSS.n968 VSS.n716 0.939203
R3092 VSS.n716 VSS.n715 0.939203
R3093 VSS.n976 VSS.n975 0.939203
R3094 VSS.n753 VSS.n740 0.939203
R3095 VSS.n744 VSS.n740 0.939203
R3096 VSS.n760 VSS.n740 0.939203
R3097 VSS.n763 VSS.n740 0.939203
R3098 VSS.n205 VSS.n200 0.939203
R3099 VSS.n1828 VSS.n247 0.939203
R3100 VSS.n1831 VSS.n247 0.939203
R3101 VSS.n1813 VSS.n247 0.939203
R3102 VSS.n1795 VSS.n247 0.939203
R3103 VSS.n1806 VSS.n247 0.939203
R3104 VSS.n1800 VSS.n247 0.939203
R3105 VSS.n2136 VSS.n169 0.939203
R3106 VSS.n2138 VSS.n169 0.939203
R3107 VSS.n2144 VSS.n169 0.939203
R3108 VSS.n2146 VSS.n169 0.939203
R3109 VSS.n2152 VSS.n169 0.939203
R3110 VSS.n2154 VSS.n169 0.939203
R3111 VSS.n2160 VSS.n169 0.939203
R3112 VSS.n2162 VSS.n169 0.939203
R3113 VSS.n2168 VSS.n169 0.939203
R3114 VSS.n2123 VSS.n169 0.939203
R3115 VSS.n2175 VSS.n169 0.939203
R3116 VSS.n1893 VSS.n47 0.939203
R3117 VSS.n1889 VSS.n47 0.939203
R3118 VSS.n2287 VSS.n47 0.939203
R3119 VSS.n2243 VSS.n47 0.939203
R3120 VSS.n2280 VSS.n47 0.939203
R3121 VSS.n2274 VSS.n47 0.939203
R3122 VSS.n2272 VSS.n2271 0.939203
R3123 VSS.n2271 VSS.n2270 0.939203
R3124 VSS.n95 VSS.n63 0.939203
R3125 VSS.n97 VSS.n63 0.939203
R3126 VSS.n103 VSS.n63 0.939203
R3127 VSS.n105 VSS.n63 0.939203
R3128 VSS.n111 VSS.n63 0.939203
R3129 VSS.n113 VSS.n63 0.939203
R3130 VSS.n119 VSS.n63 0.939203
R3131 VSS.n81 VSS.n63 0.939203
R3132 VSS.n87 VSS.n63 0.939203
R3133 VSS.n89 VSS.n63 0.939203
R3134 VSS.n227 VSS.n54 0.931463
R3135 VSS.n75 VSS.t21 0.8195
R3136 VSS.n75 VSS.t24 0.8195
R3137 VSS.n76 VSS.t20 0.8195
R3138 VSS.n76 VSS.t4 0.8195
R3139 VSS.n607 VSS.n565 0.702875
R3140 VSS.n553 VSS.n511 0.702875
R3141 VSS.n1512 VSS.n437 0.702875
R3142 VSS.n1513 VSS.n423 0.702875
R3143 VSS.n2242 VSS.n0 0.702875
R3144 VSS.n2359 VSS.n1 0.702875
R3145 VSS.n1131 VSS.n1130 0.698622
R3146 VSS.n1259 VSS.n1258 0.698622
R3147 VSS.n1387 VSS.n1386 0.698622
R3148 VSS.n1514 VSS.n436 0.698622
R3149 VSS.n1553 VSS.n341 0.698622
R3150 VSS.n2268 VSS.n43 0.698622
R3151 VSS.n2242 VSS.n2241 0.692375
R3152 VSS VSS.n607 0.629
R3153 VSS.n2241 VSS.n2240 0.624125
R3154 VSS.n565 VSS.n553 0.613625
R3155 VSS.n511 VSS.n437 0.613625
R3156 VSS.n1513 VSS.n1512 0.613625
R3157 VSS.n2359 VSS.n0 0.613625
R3158 VSS.n423 VSS.n1 0.613625
R3159 VSS.t23 VSS.n150 0.462148
R3160 VSS.n183 VSS 0.397167
R3161 VSS.n184 VSS.n183 0.367833
R3162 VSS.n1096 VSS.n1095 0.237342
R3163 VSS.n1096 VSS.n612 0.237342
R3164 VSS.n1102 VSS.n612 0.237342
R3165 VSS.n1103 VSS.n1102 0.237342
R3166 VSS.n1104 VSS.n1103 0.237342
R3167 VSS.n1104 VSS.n605 0.237342
R3168 VSS.n1124 VSS.n606 0.237342
R3169 VSS.n1124 VSS.n1123 0.237342
R3170 VSS.n1123 VSS.n1122 0.237342
R3171 VSS.n1122 VSS.n1110 0.237342
R3172 VSS.n1116 VSS.n1110 0.237342
R3173 VSS.n1116 VSS.n1115 0.237342
R3174 VSS.n1115 VSS.n1114 0.237342
R3175 VSS.n1114 VSS.n562 0.237342
R3176 VSS.n1224 VSS.n1223 0.237342
R3177 VSS.n1224 VSS.n558 0.237342
R3178 VSS.n1230 VSS.n558 0.237342
R3179 VSS.n1231 VSS.n1230 0.237342
R3180 VSS.n1232 VSS.n1231 0.237342
R3181 VSS.n1232 VSS.n551 0.237342
R3182 VSS.n1252 VSS.n552 0.237342
R3183 VSS.n1252 VSS.n1251 0.237342
R3184 VSS.n1251 VSS.n1250 0.237342
R3185 VSS.n1250 VSS.n1238 0.237342
R3186 VSS.n1244 VSS.n1238 0.237342
R3187 VSS.n1244 VSS.n1243 0.237342
R3188 VSS.n1243 VSS.n1242 0.237342
R3189 VSS.n1242 VSS.n508 0.237342
R3190 VSS.n1352 VSS.n1351 0.237342
R3191 VSS.n1352 VSS.n504 0.237342
R3192 VSS.n1358 VSS.n504 0.237342
R3193 VSS.n1359 VSS.n1358 0.237342
R3194 VSS.n1360 VSS.n1359 0.237342
R3195 VSS.n1360 VSS.n498 0.237342
R3196 VSS.n1380 VSS.n499 0.237342
R3197 VSS.n1380 VSS.n1379 0.237342
R3198 VSS.n1379 VSS.n1378 0.237342
R3199 VSS.n1378 VSS.n1366 0.237342
R3200 VSS.n1372 VSS.n1366 0.237342
R3201 VSS.n1372 VSS.n1371 0.237342
R3202 VSS.n1371 VSS.n1370 0.237342
R3203 VSS.n1370 VSS.n438 0.237342
R3204 VSS.n458 VSS.n439 0.237342
R3205 VSS.n458 VSS.n457 0.237342
R3206 VSS.n457 VSS.n456 0.237342
R3207 VSS.n456 VSS.n447 0.237342
R3208 VSS.n450 VSS.n447 0.237342
R3209 VSS.n450 VSS.n435 0.237342
R3210 VSS.n1520 VSS.n431 0.237342
R3211 VSS.n1521 VSS.n1520 0.237342
R3212 VSS.n1522 VSS.n1521 0.237342
R3213 VSS.n1522 VSS.n427 0.237342
R3214 VSS.n1529 VSS.n427 0.237342
R3215 VSS.n1530 VSS.n1529 0.237342
R3216 VSS.n1531 VSS.n1530 0.237342
R3217 VSS.n1531 VSS.n369 0.237342
R3218 VSS.n1543 VSS.n365 0.237342
R3219 VSS.n1544 VSS.n1543 0.237342
R3220 VSS.n1545 VSS.n1544 0.237342
R3221 VSS.n1545 VSS.n361 0.237342
R3222 VSS.n1551 VSS.n361 0.237342
R3223 VSS.n1552 VSS.n1551 0.237342
R3224 VSS.n1559 VSS.n357 0.237342
R3225 VSS.n1560 VSS.n1559 0.237342
R3226 VSS.n1561 VSS.n1560 0.237342
R3227 VSS.n1561 VSS.n353 0.237342
R3228 VSS.n1567 VSS.n353 0.237342
R3229 VSS.n1568 VSS.n1567 0.237342
R3230 VSS.n1569 VSS.n1568 0.237342
R3231 VSS.n1569 VSS.n2 0.237342
R3232 VSS.n2257 VSS.n3 0.237342
R3233 VSS.n2258 VSS.n2257 0.237342
R3234 VSS.n2259 VSS.n2258 0.237342
R3235 VSS.n2259 VSS.n2249 0.237342
R3236 VSS.n2265 VSS.n2249 0.237342
R3237 VSS.n2266 VSS.n2265 0.237342
R3238 VSS.n2267 VSS.n2246 0.237342
R3239 VSS.n2276 VSS.n2246 0.237342
R3240 VSS.n2277 VSS.n2276 0.237342
R3241 VSS.n2278 VSS.n2277 0.237342
R3242 VSS.n2278 VSS.n2244 0.237342
R3243 VSS.n2283 VSS.n2244 0.237342
R3244 VSS.n2284 VSS.n2283 0.237342
R3245 VSS.n2284 VSS.n51 0.237342
R3246 VSS.n1891 VSS.n52 0.237342
R3247 VSS.n1891 VSS.n1888 0.237342
R3248 VSS.n1896 VSS.n1888 0.237342
R3249 VSS.n1898 VSS.n1896 0.237342
R3250 VSS.n1899 VSS.n1898 0.237342
R3251 VSS.n1901 VSS.n1899 0.237342
R3252 VSS.n1901 VSS.n1900 0.237342
R3253 VSS.n1918 VSS.n226 0.237342
R3254 VSS.n1919 VSS.n1918 0.237342
R3255 VSS.n1938 VSS.n1919 0.237342
R3256 VSS.n1938 VSS.n1937 0.237342
R3257 VSS.n1937 VSS.n1936 0.237342
R3258 VSS.n1936 VSS.n1920 0.237342
R3259 VSS.n1920 VSS.n56 0.237342
R3260 VSS.n129 VSS.n57 0.237342
R3261 VSS.n139 VSS.n129 0.237342
R3262 VSS.n140 VSS.n139 0.237342
R3263 VSS.n2216 VSS.n140 0.237342
R3264 VSS.n2216 VSS.n2215 0.237342
R3265 VSS.n2215 VSS.n2214 0.237342
R3266 VSS.n2214 VSS.n141 0.237342
R3267 VSS.n144 VSS.n141 0.237342
R3268 VSS.n154 VSS.n144 0.237342
R3269 VSS.n155 VSS.n154 0.237342
R3270 VSS.n2199 VSS.n155 0.237342
R3271 VSS.n2199 VSS.n2198 0.237342
R3272 VSS.n2198 VSS.n2197 0.237342
R3273 VSS.n2197 VSS.n156 0.237342
R3274 VSS.n2184 VSS.n156 0.237342
R3275 VSS.n2185 VSS.n2184 0.237342
R3276 VSS.n2158 VSS.n2126 0.237342
R3277 VSS.n2158 VSS.n2157 0.237342
R3278 VSS.n2157 VSS.n2156 0.237342
R3279 VSS.n2156 VSS.n2130 0.237342
R3280 VSS.n2150 VSS.n2130 0.237342
R3281 VSS.n2148 VSS.n2132 0.237342
R3282 VSS.n2142 VSS.n2132 0.237342
R3283 VSS.n2142 VSS.n2141 0.237342
R3284 VSS.n2141 VSS.n2140 0.237342
R3285 VSS.n2140 VSS.n2135 0.237342
R3286 VSS.n2135 VSS.n2134 0.237342
R3287 VSS.n741 VSS.n721 0.237342
R3288 VSS.n758 VSS.n741 0.237342
R3289 VSS.n758 VSS.n757 0.237342
R3290 VSS.n757 VSS.n756 0.237342
R3291 VSS.n756 VSS.n743 0.237342
R3292 VSS.n751 VSS.n743 0.237342
R3293 VSS.n751 VSS.n750 0.237342
R3294 VSS.n750 VSS.n749 0.237342
R3295 VSS.n749 VSS.n689 0.237342
R3296 VSS.n1041 VSS.n689 0.237342
R3297 VSS.n1041 VSS.n1040 0.237342
R3298 VSS.n1040 VSS.n1039 0.237342
R3299 VSS.n1039 VSS.n690 0.237342
R3300 VSS.n1033 VSS.n690 0.237342
R3301 VSS.n1033 VSS.n1032 0.237342
R3302 VSS.n1032 VSS.n1031 0.237342
R3303 VSS.n122 VSS.n67 0.237342
R3304 VSS.n117 VSS.n67 0.237342
R3305 VSS.n117 VSS.n116 0.237342
R3306 VSS.n116 VSS.n115 0.237342
R3307 VSS.n115 VSS.n69 0.237342
R3308 VSS.n109 VSS.n69 0.237342
R3309 VSS.n109 VSS.n108 0.237342
R3310 VSS.n108 VSS.n107 0.237342
R3311 VSS.n107 VSS.n71 0.237342
R3312 VSS.n101 VSS.n71 0.237342
R3313 VSS.n101 VSS.n100 0.237342
R3314 VSS.n100 VSS.n99 0.237342
R3315 VSS.n99 VSS.n73 0.237342
R3316 VSS.n988 VSS.n706 0.237342
R3317 VSS.n988 VSS.n987 0.237342
R3318 VSS.n987 VSS.n986 0.237342
R3319 VSS.n986 VSS.n707 0.237342
R3320 VSS.n980 VSS.n707 0.237342
R3321 VSS.n980 VSS.n979 0.237342
R3322 VSS.n979 VSS.n978 0.237342
R3323 VSS.n978 VSS.n711 0.237342
R3324 VSS.n973 VSS.n711 0.237342
R3325 VSS.n973 VSS.n972 0.237342
R3326 VSS.n972 VSS.n971 0.237342
R3327 VSS.n971 VSS.n714 0.237342
R3328 VSS.n966 VSS.n714 0.237342
R3329 VSS.n966 VSS.n965 0.237342
R3330 VSS.n965 VSS.n964 0.237342
R3331 VSS.n964 VSS.n718 0.237342
R3332 VSS.n2087 VSS.n2085 0.237342
R3333 VSS.n2087 VSS.n2086 0.237342
R3334 VSS.n2086 VSS.n178 0.237342
R3335 VSS.n2094 VSS.n178 0.237342
R3336 VSS.n2095 VSS.n2094 0.237342
R3337 VSS.n2095 VSS.n176 0.237342
R3338 VSS.n2100 VSS.n176 0.237342
R3339 VSS.n2045 VSS.n2042 0.237342
R3340 VSS.n2042 VSS.n2041 0.237342
R3341 VSS.n2041 VSS.n2038 0.237342
R3342 VSS.n2038 VSS.n2037 0.237342
R3343 VSS.n2037 VSS.n2031 0.237342
R3344 VSS.n2032 VSS.n2031 0.237342
R3345 VSS.n2032 VSS.n194 0.237342
R3346 VSS.n2064 VSS.n194 0.237342
R3347 VSS.n2065 VSS.n2064 0.237342
R3348 VSS.n2066 VSS.n2065 0.237342
R3349 VSS.n2066 VSS.n190 0.237342
R3350 VSS.n2072 VSS.n190 0.237342
R3351 VSS.n2073 VSS.n2072 0.237342
R3352 VSS.n2074 VSS.n2073 0.237342
R3353 VSS.n2074 VSS.n186 0.237342
R3354 VSS.n2083 VSS.n186 0.237342
R3355 VSS.n1988 VSS.n1985 0.237342
R3356 VSS.n2025 VSS.n1988 0.237342
R3357 VSS.n2025 VSS.n2024 0.237342
R3358 VSS.n2024 VSS.n2023 0.237342
R3359 VSS.n2023 VSS.n1989 0.237342
R3360 VSS.n2017 VSS.n1989 0.237342
R3361 VSS.n2017 VSS.n2016 0.237342
R3362 VSS.n2016 VSS.n2015 0.237342
R3363 VSS.n2015 VSS.n1993 0.237342
R3364 VSS.n2008 VSS.n1993 0.237342
R3365 VSS.n2008 VSS.n2007 0.237342
R3366 VSS.n2007 VSS.n2006 0.237342
R3367 VSS.n2006 VSS.n1995 0.237342
R3368 VSS.n2001 VSS.n1995 0.237342
R3369 VSS.n2001 VSS.n2000 0.237342
R3370 VSS.n2000 VSS.n123 0.237342
R3371 VSS.n219 VSS.n216 0.237342
R3372 VSS.n1974 VSS.n219 0.237342
R3373 VSS.n1974 VSS.n1973 0.237342
R3374 VSS.n1973 VSS.n1972 0.237342
R3375 VSS.n1972 VSS.n221 0.237342
R3376 VSS.n1967 VSS.n221 0.237342
R3377 VSS.n1967 VSS.n1966 0.237342
R3378 VSS.n1966 VSS.n1965 0.237342
R3379 VSS.n1965 VSS.n1955 0.237342
R3380 VSS.n1960 VSS.n1955 0.237342
R3381 VSS.n1960 VSS.n1959 0.237342
R3382 VSS.n1959 VSS.n215 0.237342
R3383 VSS.n2058 VSS.n215 0.237342
R3384 VSS.n2058 VSS.n2057 0.237342
R3385 VSS.n2057 VSS.n2056 0.237342
R3386 VSS.n2056 VSS.n2053 0.237342
R3387 VSS.n1761 VSS.n1760 0.237342
R3388 VSS.n1762 VSS.n1761 0.237342
R3389 VSS.n1762 VSS.n262 0.237342
R3390 VSS.n1768 VSS.n262 0.237342
R3391 VSS.n1769 VSS.n1768 0.237342
R3392 VSS.n1770 VSS.n1769 0.237342
R3393 VSS.n1770 VSS.n257 0.237342
R3394 VSS.n1777 VSS.n257 0.237342
R3395 VSS.n1778 VSS.n1777 0.237342
R3396 VSS.n1779 VSS.n1778 0.237342
R3397 VSS.n1779 VSS.n253 0.237342
R3398 VSS.n1785 VSS.n253 0.237342
R3399 VSS.n1786 VSS.n1785 0.237342
R3400 VSS.n1787 VSS.n1786 0.237342
R3401 VSS.n1787 VSS.n249 0.237342
R3402 VSS.n1793 VSS.n249 0.237342
R3403 VSS.n1681 VSS.n1678 0.237342
R3404 VSS.n1678 VSS.n1677 0.237342
R3405 VSS.n1677 VSS.n1674 0.237342
R3406 VSS.n1674 VSS.n273 0.237342
R3407 VSS.n1732 VSS.n273 0.237342
R3408 VSS.n1733 VSS.n1732 0.237342
R3409 VSS.n1735 VSS.n1733 0.237342
R3410 VSS.n1735 VSS.n1734 0.237342
R3411 VSS.n1734 VSS.n270 0.237342
R3412 VSS.n1742 VSS.n270 0.237342
R3413 VSS.n1743 VSS.n1742 0.237342
R3414 VSS.n1744 VSS.n1743 0.237342
R3415 VSS.n1744 VSS.n268 0.237342
R3416 VSS.n1750 VSS.n268 0.237342
R3417 VSS.n1751 VSS.n1750 0.237342
R3418 VSS.n1752 VSS.n1751 0.237342
R3419 VSS.n1726 VSS.n1725 0.237342
R3420 VSS.n1725 VSS.n1724 0.237342
R3421 VSS.n1724 VSS.n1686 0.237342
R3422 VSS.n1718 VSS.n1686 0.237342
R3423 VSS.n1718 VSS.n1717 0.237342
R3424 VSS.n1717 VSS.n1716 0.237342
R3425 VSS.n1716 VSS.n1690 0.237342
R3426 VSS.n1692 VSS.n1690 0.237342
R3427 VSS.n1695 VSS.n1692 0.237342
R3428 VSS.n1706 VSS.n1695 0.237342
R3429 VSS.n1706 VSS.n1705 0.237342
R3430 VSS.n1705 VSS.n1704 0.237342
R3431 VSS.n1704 VSS.n1700 0.237342
R3432 VSS.n1700 VSS.n1699 0.237342
R3433 VSS.n1699 VSS.n1696 0.237342
R3434 VSS.n1696 VSS.n31 0.237342
R3435 VSS.n301 VSS.n298 0.237342
R3436 VSS.n302 VSS.n301 0.237342
R3437 VSS.n303 VSS.n302 0.237342
R3438 VSS.n303 VSS.n289 0.237342
R3439 VSS.n1649 VSS.n289 0.237342
R3440 VSS.n1650 VSS.n1649 0.237342
R3441 VSS.n1652 VSS.n1650 0.237342
R3442 VSS.n1652 VSS.n1651 0.237342
R3443 VSS.n1651 VSS.n286 0.237342
R3444 VSS.n1658 VSS.n286 0.237342
R3445 VSS.n1659 VSS.n1658 0.237342
R3446 VSS.n1662 VSS.n1659 0.237342
R3447 VSS.n1663 VSS.n1662 0.237342
R3448 VSS.n1666 VSS.n1663 0.237342
R3449 VSS.n1667 VSS.n1666 0.237342
R3450 VSS.n1670 VSS.n1667 0.237342
R3451 VSS.n1643 VSS.n1642 0.237342
R3452 VSS.n1642 VSS.n1641 0.237342
R3453 VSS.n1641 VSS.n312 0.237342
R3454 VSS.n1635 VSS.n312 0.237342
R3455 VSS.n1635 VSS.n1634 0.237342
R3456 VSS.n1634 VSS.n1633 0.237342
R3457 VSS.n1633 VSS.n316 0.237342
R3458 VSS.n1626 VSS.n316 0.237342
R3459 VSS.n1626 VSS.n1625 0.237342
R3460 VSS.n1625 VSS.n1624 0.237342
R3461 VSS.n1624 VSS.n321 0.237342
R3462 VSS.n1618 VSS.n321 0.237342
R3463 VSS.n1618 VSS.n1617 0.237342
R3464 VSS.n1617 VSS.n1616 0.237342
R3465 VSS.n1616 VSS.n325 0.237342
R3466 VSS.n1611 VSS.n325 0.237342
R3467 VSS.n918 VSS.n917 0.237342
R3468 VSS.n917 VSS.n916 0.237342
R3469 VSS.n916 VSS.n879 0.237342
R3470 VSS.n911 VSS.n879 0.237342
R3471 VSS.n911 VSS.n910 0.237342
R3472 VSS.n910 VSS.n909 0.237342
R3473 VSS.n909 VSS.n882 0.237342
R3474 VSS.n886 VSS.n882 0.237342
R3475 VSS.n903 VSS.n886 0.237342
R3476 VSS.n903 VSS.n902 0.237342
R3477 VSS.n902 VSS.n901 0.237342
R3478 VSS.n901 VSS.n898 0.237342
R3479 VSS.n898 VSS.n897 0.237342
R3480 VSS.n897 VSS.n894 0.237342
R3481 VSS.n894 VSS.n893 0.237342
R3482 VSS.n893 VSS.n890 0.237342
R3483 VSS.n876 VSS.n832 0.237342
R3484 VSS.n870 VSS.n832 0.237342
R3485 VSS.n870 VSS.n869 0.237342
R3486 VSS.n869 VSS.n868 0.237342
R3487 VSS.n868 VSS.n836 0.237342
R3488 VSS.n862 VSS.n836 0.237342
R3489 VSS.n862 VSS.n861 0.237342
R3490 VSS.n861 VSS.n860 0.237342
R3491 VSS.n860 VSS.n840 0.237342
R3492 VSS.n854 VSS.n840 0.237342
R3493 VSS.n854 VSS.n853 0.237342
R3494 VSS.n853 VSS.n852 0.237342
R3495 VSS.n852 VSS.n848 0.237342
R3496 VSS.n848 VSS.n847 0.237342
R3497 VSS.n847 VSS.n844 0.237342
R3498 VSS.n844 VSS.n484 0.237342
R3499 VSS.n953 VSS.n952 0.237342
R3500 VSS.n952 VSS.n951 0.237342
R3501 VSS.n951 VSS.n816 0.237342
R3502 VSS.n946 VSS.n816 0.237342
R3503 VSS.n946 VSS.n945 0.237342
R3504 VSS.n945 VSS.n944 0.237342
R3505 VSS.n944 VSS.n819 0.237342
R3506 VSS.n823 VSS.n819 0.237342
R3507 VSS.n938 VSS.n823 0.237342
R3508 VSS.n938 VSS.n937 0.237342
R3509 VSS.n937 VSS.n936 0.237342
R3510 VSS.n936 VSS.n824 0.237342
R3511 VSS.n931 VSS.n824 0.237342
R3512 VSS.n931 VSS.n930 0.237342
R3513 VSS.n930 VSS.n929 0.237342
R3514 VSS.n929 VSS.n828 0.237342
R3515 VSS.n813 VSS.n768 0.237342
R3516 VSS.n807 VSS.n768 0.237342
R3517 VSS.n807 VSS.n806 0.237342
R3518 VSS.n806 VSS.n805 0.237342
R3519 VSS.n805 VSS.n772 0.237342
R3520 VSS.n799 VSS.n772 0.237342
R3521 VSS.n799 VSS.n798 0.237342
R3522 VSS.n798 VSS.n797 0.237342
R3523 VSS.n797 VSS.n776 0.237342
R3524 VSS.n791 VSS.n776 0.237342
R3525 VSS.n791 VSS.n790 0.237342
R3526 VSS.n790 VSS.n789 0.237342
R3527 VSS.n789 VSS.n785 0.237342
R3528 VSS.n785 VSS.n784 0.237342
R3529 VSS.n784 VSS.n781 0.237342
R3530 VSS.n781 VSS.n537 0.237342
R3531 VSS.n1025 VSS.n1024 0.237342
R3532 VSS.n1024 VSS.n1023 0.237342
R3533 VSS.n1023 VSS.n1020 0.237342
R3534 VSS.n1020 VSS.n1019 0.237342
R3535 VSS.n1019 VSS.n1016 0.237342
R3536 VSS.n1016 VSS.n1015 0.237342
R3537 VSS.n1015 VSS.n1012 0.237342
R3538 VSS.n1012 VSS.n1011 0.237342
R3539 VSS.n1011 VSS.n1008 0.237342
R3540 VSS.n1008 VSS.n1007 0.237342
R3541 VSS.n1007 VSS.n1004 0.237342
R3542 VSS.n1004 VSS.n1003 0.237342
R3543 VSS.n1003 VSS.n1000 0.237342
R3544 VSS.n1000 VSS.n999 0.237342
R3545 VSS.n999 VSS.n996 0.237342
R3546 VSS.n996 VSS.n591 0.237342
R3547 VSS.n674 VSS.n623 0.237342
R3548 VSS.n669 VSS.n623 0.237342
R3549 VSS.n669 VSS.n668 0.237342
R3550 VSS.n668 VSS.n625 0.237342
R3551 VSS.n663 VSS.n625 0.237342
R3552 VSS.n663 VSS.n662 0.237342
R3553 VSS.n662 VSS.n661 0.237342
R3554 VSS.n661 VSS.n627 0.237342
R3555 VSS.n655 VSS.n627 0.237342
R3556 VSS.n655 VSS.n654 0.237342
R3557 VSS.n654 VSS.n653 0.237342
R3558 VSS.n653 VSS.n629 0.237342
R3559 VSS.n647 VSS.n629 0.237342
R3560 VSS.n647 VSS.n646 0.237342
R3561 VSS.n646 VSS.n645 0.237342
R3562 VSS.n645 VSS.n631 0.237342
R3563 VSS.n640 VSS.n631 0.237342
R3564 VSS.n640 VSS.n639 0.237342
R3565 VSS.n639 VSS.n633 0.237342
R3566 VSS.n634 VSS.n633 0.237342
R3567 VSS.n634 VSS.n616 0.237342
R3568 VSS.n1205 VSS.n1204 0.237342
R3569 VSS.n1204 VSS.n1203 0.237342
R3570 VSS.n1203 VSS.n1200 0.237342
R3571 VSS.n1200 VSS.n1199 0.237342
R3572 VSS.n1199 VSS.n1196 0.237342
R3573 VSS.n1196 VSS.n1195 0.237342
R3574 VSS.n1195 VSS.n1192 0.237342
R3575 VSS.n1192 VSS.n1191 0.237342
R3576 VSS.n1191 VSS.n1188 0.237342
R3577 VSS.n1188 VSS.n1187 0.237342
R3578 VSS.n1187 VSS.n1184 0.237342
R3579 VSS.n1184 VSS.n1183 0.237342
R3580 VSS.n1183 VSS.n1180 0.237342
R3581 VSS.n1180 VSS.n575 0.237342
R3582 VSS.n1210 VSS.n575 0.237342
R3583 VSS.n1211 VSS.n1210 0.237342
R3584 VSS.n1217 VSS.n1211 0.237342
R3585 VSS.n1217 VSS.n1216 0.237342
R3586 VSS.n1216 VSS.n1215 0.237342
R3587 VSS.n1215 VSS.n1212 0.237342
R3588 VSS.n1212 VSS.n563 0.237342
R3589 VSS.n1333 VSS.n1332 0.237342
R3590 VSS.n1332 VSS.n1331 0.237342
R3591 VSS.n1331 VSS.n1328 0.237342
R3592 VSS.n1328 VSS.n1327 0.237342
R3593 VSS.n1327 VSS.n1324 0.237342
R3594 VSS.n1324 VSS.n1323 0.237342
R3595 VSS.n1323 VSS.n1320 0.237342
R3596 VSS.n1320 VSS.n1319 0.237342
R3597 VSS.n1319 VSS.n1316 0.237342
R3598 VSS.n1316 VSS.n1315 0.237342
R3599 VSS.n1315 VSS.n1312 0.237342
R3600 VSS.n1312 VSS.n1311 0.237342
R3601 VSS.n1311 VSS.n1308 0.237342
R3602 VSS.n1308 VSS.n521 0.237342
R3603 VSS.n1338 VSS.n521 0.237342
R3604 VSS.n1339 VSS.n1338 0.237342
R3605 VSS.n1345 VSS.n1339 0.237342
R3606 VSS.n1345 VSS.n1344 0.237342
R3607 VSS.n1344 VSS.n1343 0.237342
R3608 VSS.n1343 VSS.n1340 0.237342
R3609 VSS.n1340 VSS.n509 0.237342
R3610 VSS.n1494 VSS.n1493 0.237342
R3611 VSS.n1493 VSS.n1492 0.237342
R3612 VSS.n1492 VSS.n1489 0.237342
R3613 VSS.n1489 VSS.n1488 0.237342
R3614 VSS.n1488 VSS.n1485 0.237342
R3615 VSS.n1485 VSS.n1484 0.237342
R3616 VSS.n1484 VSS.n1481 0.237342
R3617 VSS.n1481 VSS.n1480 0.237342
R3618 VSS.n1480 VSS.n1477 0.237342
R3619 VSS.n1477 VSS.n1476 0.237342
R3620 VSS.n1476 VSS.n1473 0.237342
R3621 VSS.n1473 VSS.n1472 0.237342
R3622 VSS.n1472 VSS.n1469 0.237342
R3623 VSS.n1469 VSS.n468 0.237342
R3624 VSS.n1499 VSS.n468 0.237342
R3625 VSS.n1500 VSS.n1499 0.237342
R3626 VSS.n1506 VSS.n1500 0.237342
R3627 VSS.n1506 VSS.n1505 0.237342
R3628 VSS.n1505 VSS.n1504 0.237342
R3629 VSS.n1504 VSS.n1501 0.237342
R3630 VSS.n1501 VSS.n440 0.237342
R3631 VSS.n384 VSS.n329 0.237342
R3632 VSS.n385 VSS.n384 0.237342
R3633 VSS.n386 VSS.n385 0.237342
R3634 VSS.n386 VSS.n379 0.237342
R3635 VSS.n392 VSS.n379 0.237342
R3636 VSS.n393 VSS.n392 0.237342
R3637 VSS.n394 VSS.n393 0.237342
R3638 VSS.n394 VSS.n377 0.237342
R3639 VSS.n400 VSS.n377 0.237342
R3640 VSS.n401 VSS.n400 0.237342
R3641 VSS.n402 VSS.n401 0.237342
R3642 VSS.n402 VSS.n375 0.237342
R3643 VSS.n408 VSS.n375 0.237342
R3644 VSS.n409 VSS.n408 0.237342
R3645 VSS.n410 VSS.n409 0.237342
R3646 VSS.n410 VSS.n373 0.237342
R3647 VSS.n373 VSS.n372 0.237342
R3648 VSS.n416 VSS.n372 0.237342
R3649 VSS.n417 VSS.n416 0.237342
R3650 VSS.n417 VSS.n370 0.237342
R3651 VSS.n422 VSS.n370 0.237342
R3652 VSS.n1835 VSS.n245 0.237342
R3653 VSS.n1841 VSS.n245 0.237342
R3654 VSS.n1842 VSS.n1841 0.237342
R3655 VSS.n1843 VSS.n1842 0.237342
R3656 VSS.n1843 VSS.n240 0.237342
R3657 VSS.n1850 VSS.n240 0.237342
R3658 VSS.n1851 VSS.n1850 0.237342
R3659 VSS.n1883 VSS.n1851 0.237342
R3660 VSS.n1883 VSS.n1882 0.237342
R3661 VSS.n1882 VSS.n1881 0.237342
R3662 VSS.n1881 VSS.n1852 0.237342
R3663 VSS.n1875 VSS.n1852 0.237342
R3664 VSS.n1875 VSS.n1874 0.237342
R3665 VSS.n1874 VSS.n1873 0.237342
R3666 VSS.n1873 VSS.n1856 0.237342
R3667 VSS.n1867 VSS.n1856 0.237342
R3668 VSS.n1867 VSS.n1866 0.237342
R3669 VSS.n1866 VSS.n1865 0.237342
R3670 VSS.n1865 VSS.n1860 0.237342
R3671 VSS.n1860 VSS.n50 0.237342
R3672 VSS.n2290 VSS.n50 0.237342
R3673 VSS.n2341 VSS.n2340 0.237342
R3674 VSS.n2340 VSS.n2339 0.237342
R3675 VSS.n2339 VSS.n2336 0.237342
R3676 VSS.n2336 VSS.n2335 0.237342
R3677 VSS.n2335 VSS.n2332 0.237342
R3678 VSS.n2332 VSS.n2331 0.237342
R3679 VSS.n2331 VSS.n2328 0.237342
R3680 VSS.n2328 VSS.n2327 0.237342
R3681 VSS.n2327 VSS.n2324 0.237342
R3682 VSS.n2324 VSS.n2323 0.237342
R3683 VSS.n2323 VSS.n2320 0.237342
R3684 VSS.n2320 VSS.n2319 0.237342
R3685 VSS.n2319 VSS.n2316 0.237342
R3686 VSS.n2316 VSS.n15 0.237342
R3687 VSS.n2346 VSS.n15 0.237342
R3688 VSS.n2347 VSS.n2346 0.237342
R3689 VSS.n2353 VSS.n2347 0.237342
R3690 VSS.n2353 VSS.n2352 0.237342
R3691 VSS.n2352 VSS.n2351 0.237342
R3692 VSS.n2351 VSS.n2348 0.237342
R3693 VSS.n2348 VSS.n4 0.237342
R3694 VSS.n2106 VSS.n2105 0.237342
R3695 VSS.n2106 VSS.n174 0.237342
R3696 VSS.n2112 VSS.n174 0.237342
R3697 VSS.n2113 VSS.n2112 0.237342
R3698 VSS.n2114 VSS.n2113 0.237342
R3699 VSS.n2114 VSS.n172 0.237342
R3700 VSS.n172 VSS.n171 0.237342
R3701 VSS.n2121 VSS.n171 0.237342
R3702 VSS.n2177 VSS.n2122 0.237342
R3703 VSS.n2172 VSS.n2122 0.237342
R3704 VSS.n2172 VSS.n2171 0.237342
R3705 VSS.n2171 VSS.n2124 0.237342
R3706 VSS.n2166 VSS.n2124 0.237342
R3707 VSS.n2166 VSS.n2165 0.237342
R3708 VSS.n1088 VSS.n1087 0.237342
R3709 VSS.n1087 VSS.n1086 0.237342
R3710 VSS.n1086 VSS.n1068 0.237342
R3711 VSS.n1080 VSS.n1068 0.237342
R3712 VSS.n1080 VSS.n1079 0.237342
R3713 VSS.n1079 VSS.n1078 0.237342
R3714 VSS.n1078 VSS.n1073 0.237342
R3715 VSS.n1073 VSS.n602 0.237342
R3716 VSS.n1135 VSS.n602 0.237342
R3717 VSS.n1136 VSS.n1135 0.237342
R3718 VSS.n1137 VSS.n1136 0.237342
R3719 VSS.n1137 VSS.n598 0.237342
R3720 VSS.n1143 VSS.n598 0.237342
R3721 VSS.n1144 VSS.n1143 0.237342
R3722 VSS.n1146 VSS.n1144 0.237342
R3723 VSS.n1146 VSS.n1145 0.237342
R3724 VSS.n1145 VSS.n592 0.237342
R3725 VSS.n1154 VSS.n592 0.237342
R3726 VSS.n1178 VSS.n1155 0.237342
R3727 VSS.n1172 VSS.n1155 0.237342
R3728 VSS.n1172 VSS.n1171 0.237342
R3729 VSS.n1171 VSS.n1170 0.237342
R3730 VSS.n1170 VSS.n1159 0.237342
R3731 VSS.n1164 VSS.n1159 0.237342
R3732 VSS.n1164 VSS.n1163 0.237342
R3733 VSS.n1163 VSS.n548 0.237342
R3734 VSS.n1263 VSS.n548 0.237342
R3735 VSS.n1264 VSS.n1263 0.237342
R3736 VSS.n1265 VSS.n1264 0.237342
R3737 VSS.n1265 VSS.n544 0.237342
R3738 VSS.n1271 VSS.n544 0.237342
R3739 VSS.n1272 VSS.n1271 0.237342
R3740 VSS.n1274 VSS.n1272 0.237342
R3741 VSS.n1274 VSS.n1273 0.237342
R3742 VSS.n1273 VSS.n538 0.237342
R3743 VSS.n1282 VSS.n538 0.237342
R3744 VSS.n1306 VSS.n1283 0.237342
R3745 VSS.n1300 VSS.n1283 0.237342
R3746 VSS.n1300 VSS.n1299 0.237342
R3747 VSS.n1299 VSS.n1298 0.237342
R3748 VSS.n1298 VSS.n1287 0.237342
R3749 VSS.n1292 VSS.n1287 0.237342
R3750 VSS.n1292 VSS.n1291 0.237342
R3751 VSS.n1291 VSS.n495 0.237342
R3752 VSS.n1391 VSS.n495 0.237342
R3753 VSS.n1392 VSS.n1391 0.237342
R3754 VSS.n1393 VSS.n1392 0.237342
R3755 VSS.n1393 VSS.n491 0.237342
R3756 VSS.n1399 VSS.n491 0.237342
R3757 VSS.n1400 VSS.n1399 0.237342
R3758 VSS.n1402 VSS.n1400 0.237342
R3759 VSS.n1402 VSS.n1401 0.237342
R3760 VSS.n1401 VSS.n485 0.237342
R3761 VSS.n1410 VSS.n485 0.237342
R3762 VSS.n1467 VSS.n1411 0.237342
R3763 VSS.n1461 VSS.n1411 0.237342
R3764 VSS.n1461 VSS.n1460 0.237342
R3765 VSS.n1460 VSS.n1459 0.237342
R3766 VSS.n1459 VSS.n1415 0.237342
R3767 VSS.n1453 VSS.n1415 0.237342
R3768 VSS.n1453 VSS.n1452 0.237342
R3769 VSS.n1452 VSS.n1451 0.237342
R3770 VSS.n1451 VSS.n1419 0.237342
R3771 VSS.n1444 VSS.n1419 0.237342
R3772 VSS.n1444 VSS.n1443 0.237342
R3773 VSS.n1443 VSS.n1442 0.237342
R3774 VSS.n1442 VSS.n1423 0.237342
R3775 VSS.n1436 VSS.n1423 0.237342
R3776 VSS.n1436 VSS.n1435 0.237342
R3777 VSS.n1435 VSS.n1434 0.237342
R3778 VSS.n1434 VSS.n1427 0.237342
R3779 VSS.n1427 VSS.n330 0.237342
R3780 VSS.n1609 VSS.n331 0.237342
R3781 VSS.n1603 VSS.n331 0.237342
R3782 VSS.n1603 VSS.n1602 0.237342
R3783 VSS.n1602 VSS.n1601 0.237342
R3784 VSS.n1601 VSS.n335 0.237342
R3785 VSS.n1595 VSS.n335 0.237342
R3786 VSS.n1595 VSS.n1594 0.237342
R3787 VSS.n1594 VSS.n1593 0.237342
R3788 VSS.n1593 VSS.n339 0.237342
R3789 VSS.n1586 VSS.n339 0.237342
R3790 VSS.n1586 VSS.n1585 0.237342
R3791 VSS.n1585 VSS.n1584 0.237342
R3792 VSS.n1584 VSS.n344 0.237342
R3793 VSS.n1578 VSS.n344 0.237342
R3794 VSS.n1578 VSS.n1577 0.237342
R3795 VSS.n1577 VSS.n1576 0.237342
R3796 VSS.n1576 VSS.n348 0.237342
R3797 VSS.n348 VSS.n32 0.237342
R3798 VSS.n2314 VSS.n33 0.237342
R3799 VSS.n2308 VSS.n33 0.237342
R3800 VSS.n2308 VSS.n2307 0.237342
R3801 VSS.n2307 VSS.n2306 0.237342
R3802 VSS.n2306 VSS.n37 0.237342
R3803 VSS.n2300 VSS.n37 0.237342
R3804 VSS.n2300 VSS.n2299 0.237342
R3805 VSS.n2299 VSS.n2298 0.237342
R3806 VSS.n2298 VSS.n41 0.237342
R3807 VSS.n1798 VSS.n41 0.237342
R3808 VSS.n1802 VSS.n1798 0.237342
R3809 VSS.n1803 VSS.n1802 0.237342
R3810 VSS.n1804 VSS.n1803 0.237342
R3811 VSS.n1804 VSS.n1796 0.237342
R3812 VSS.n1809 VSS.n1796 0.237342
R3813 VSS.n1810 VSS.n1809 0.237342
R3814 VSS.n1810 VSS.n1794 0.237342
R3815 VSS.n1815 VSS.n1794 0.237342
R3816 VSS.n1833 VSS.n1816 0.237342
R3817 VSS.n1817 VSS.n1816 0.237342
R3818 VSS.n1826 VSS.n1817 0.237342
R3819 VSS.n1826 VSS.n1825 0.237342
R3820 VSS.n1825 VSS.n1824 0.237342
R3821 VSS.n1824 VSS.n1819 0.237342
R3822 VSS.n1819 VSS.n232 0.237342
R3823 VSS.n1909 VSS.n232 0.237342
R3824 VSS.n1910 VSS.n1909 0.237342
R3825 VSS.n1945 VSS.n1910 0.237342
R3826 VSS.n1945 VSS.n1944 0.237342
R3827 VSS.n1944 VSS.n1943 0.237342
R3828 VSS.n1943 VSS.n1911 0.237342
R3829 VSS.n1929 VSS.n1911 0.237342
R3830 VSS.n1931 VSS.n1929 0.237342
R3831 VSS.n1931 VSS.n1930 0.237342
R3832 VSS.n1930 VSS.n66 0.237342
R3833 VSS.n2234 VSS.n66 0.237342
R3834 VSS.n2232 VSS.n124 0.237342
R3835 VSS.n2223 VSS.n124 0.237342
R3836 VSS.n2223 VSS.n2222 0.237342
R3837 VSS.n2222 VSS.n2221 0.237342
R3838 VSS.n2221 VSS.n132 0.237342
R3839 VSS.n203 VSS.n132 0.237342
R3840 VSS.n203 VSS.n202 0.237342
R3841 VSS.n202 VSS.n147 0.237342
R3842 VSS.n2206 VSS.n147 0.237342
R3843 VSS.n2206 VSS.n2205 0.237342
R3844 VSS.n2205 VSS.n2204 0.237342
R3845 VSS.n2204 VSS.n148 0.237342
R3846 VSS.n162 VSS.n148 0.237342
R3847 VSS.n2192 VSS.n162 0.237342
R3848 VSS.n2192 VSS.n2191 0.237342
R3849 VSS.n2191 VSS.n2190 0.237342
R3850 VSS.n2190 VSS.n163 0.237342
R3851 VSS.n2179 VSS.n163 0.237342
R3852 VSS.n736 VSS.n722 0.237342
R3853 VSS.n736 VSS.n735 0.237342
R3854 VSS.n735 VSS.n734 0.237342
R3855 VSS.n734 VSS.n726 0.237342
R3856 VSS.n728 VSS.n726 0.237342
R3857 VSS.n728 VSS.n682 0.237342
R3858 VSS.n1048 VSS.n682 0.237342
R3859 VSS.n1049 VSS.n1048 0.237342
R3860 VSS.n1050 VSS.n1049 0.237342
R3861 VSS.n1050 VSS.n678 0.237342
R3862 VSS.n1057 VSS.n678 0.237342
R3863 VSS.n1058 VSS.n1057 0.237342
R3864 VSS.n1059 VSS.n1058 0.237342
R3865 VSS.n1059 VSS.n676 0.237342
R3866 VSS.n676 VSS.n675 0.237342
R3867 VSS.n1066 VSS.n675 0.237342
R3868 VSS.n92 VSS.n91 0.237342
R3869 VSS.n91 VSS.n78 0.237342
R3870 VSS.n85 VSS.n78 0.237342
R3871 VSS.n85 VSS.n84 0.237342
R3872 VSS.n84 VSS.n83 0.237342
R3873 VSS.n83 VSS.n58 0.237342
R3874 VSS.n1130 VSS.n605 0.216026
R3875 VSS.n1258 VSS.n551 0.216026
R3876 VSS.n1386 VSS.n498 0.216026
R3877 VSS.n1514 VSS.n435 0.216026
R3878 VSS.n1553 VSS.n1552 0.216026
R3879 VSS.n2268 VSS.n2266 0.216026
R3880 VSS.n1900 VSS.n54 0.206553
R3881 VSS.n1095 VSS.n1094 0.192342
R3882 VSS.n1223 VSS.n1222 0.192342
R3883 VSS.n1351 VSS.n1350 0.192342
R3884 VSS.n1511 VSS.n439 0.192342
R3885 VSS.n1537 VSS.n365 0.192342
R3886 VSS.n2358 VSS.n3 0.192342
R3887 VSS.n2289 VSS.n52 0.192342
R3888 VSS.n2239 VSS.n57 0.192342
R3889 VSS.n765 VSS.n721 0.192342
R3890 VSS.n706 VSS.n694 0.192342
R3891 VSS.n2046 VSS.n2045 0.192342
R3892 VSS.n1982 VSS.n216 0.192342
R3893 VSS.n1682 VSS.n1681 0.192342
R3894 VSS.n298 VSS.n285 0.192342
R3895 VSS.n918 VSS.n877 0.192342
R3896 VSS.n953 VSS.n814 0.192342
R3897 VSS.n1222 VSS.n562 0.173395
R3898 VSS.n1350 VSS.n508 0.173395
R3899 VSS.n1511 VSS.n438 0.173395
R3900 VSS.n1537 VSS.n369 0.173395
R3901 VSS.n2358 VSS.n2 0.173395
R3902 VSS.n2289 VSS.n51 0.173395
R3903 VSS.n2239 VSS.n56 0.173395
R3904 VSS.n2185 VSS.n55 0.173395
R3905 VSS.n1031 VSS.n694 0.173395
R3906 VSS.n767 VSS.n718 0.173395
R3907 VSS.n2084 VSS.n2083 0.173395
R3908 VSS.n2053 VSS.n2052 0.173395
R3909 VSS.n1752 VSS.n266 0.173395
R3910 VSS.n1671 VSS.n1670 0.173395
R3911 VSS.n890 VSS.n889 0.173395
R3912 VSS.n831 VSS.n828 0.173395
R3913 VSS.n93 VSS.n73 0.161553
R3914 VSS.n1088 VSS.n1067 0.161553
R3915 VSS.n1179 VSS.n1178 0.161553
R3916 VSS.n1307 VSS.n1306 0.161553
R3917 VSS.n1468 VSS.n1467 0.161553
R3918 VSS.n1610 VSS.n1609 0.161553
R3919 VSS.n2315 VSS.n2314 0.161553
R3920 VSS.n1834 VSS.n1833 0.161553
R3921 VSS.n2233 VSS.n2232 0.161553
R3922 VSS.n2150 VSS.n2149 0.137868
R3923 VSS.n1094 VSS 0.124325
R3924 VSS.n2134 VSS.n55 0.119442
R3925 VSS.n1094 VSS.n616 0.119442
R3926 VSS.n1179 VSS.n1154 0.114184
R3927 VSS.n1307 VSS.n1282 0.114184
R3928 VSS.n1468 VSS.n1410 0.114184
R3929 VSS.n1610 VSS.n330 0.114184
R3930 VSS.n2315 VSS.n32 0.114184
R3931 VSS.n1834 VSS.n1815 0.114184
R3932 VSS.n2234 VSS.n2233 0.114184
R3933 VSS.n2179 VSS.n2178 0.114184
R3934 VSS.n2105 VSS.n2104 0.113
R3935 VSS.n1222 VSS.n563 0.112898
R3936 VSS.n1350 VSS.n509 0.112898
R3937 VSS.n1511 VSS.n440 0.112898
R3938 VSS.n1537 VSS.n422 0.112898
R3939 VSS.n2290 VSS.n2289 0.112898
R3940 VSS.n2358 VSS.n4 0.112898
R3941 VSS.n2239 VSS.n58 0.112898
R3942 VSS.n1130 VSS.n607 0.112876
R3943 VSS.n1258 VSS.n553 0.112876
R3944 VSS.n1386 VSS.n437 0.112876
R3945 VSS.n1514 VSS.n1513 0.112876
R3946 VSS.n1553 VSS.n1 0.112876
R3947 VSS.n2268 VSS.n0 0.112876
R3948 VSS.n2233 VSS.n122 0.101158
R3949 VSS.n1067 VSS.n674 0.101158
R3950 VSS.n1205 VSS.n1179 0.101158
R3951 VSS.n1333 VSS.n1307 0.101158
R3952 VSS.n1494 VSS.n1468 0.101158
R3953 VSS.n1610 VSS.n329 0.101158
R3954 VSS.n1835 VSS.n1834 0.101158
R3955 VSS.n2341 VSS.n2315 0.101158
R3956 VSS.n2178 VSS.n2177 0.101158
R3957 VSS.n765 VSS.n722 0.100495
R3958 VSS.n2085 VSS.n2084 0.100495
R3959 VSS.n1222 VSS.n565 0.0966111
R3960 VSS.n1350 VSS.n511 0.0966111
R3961 VSS.n1512 VSS.n1511 0.0966111
R3962 VSS.n1537 VSS.n423 0.0966111
R3963 VSS.n2289 VSS.n2242 0.0966111
R3964 VSS.n2359 VSS.n2358 0.0966111
R3965 VSS.n2240 VSS.n2239 0.0966111
R3966 VSS.n1025 VSS.n694 0.0939503
R3967 VSS.n2241 VSS.n54 0.0938027
R3968 VSS.n2084 VSS.n184 0.093725
R3969 VSS VSS.n765 0.089225
R3970 VSS.n1985 VSS.n1983 0.0833947
R3971 VSS.n1760 VSS.n1757 0.0833947
R3972 VSS.n1726 VSS.n1685 0.0833947
R3973 VSS.n1643 VSS.n311 0.0833947
R3974 VSS.n923 VSS.n876 0.0833947
R3975 VSS.n958 VSS.n813 0.0833947
R3976 VSS.n2165 VSS.n2164 0.0798421
R3977 VSS.n2164 VSS.n2126 0.0632632
R3978 VSS.n2233 VSS.n123 0.0466842
R3979 VSS.n1834 VSS.n1793 0.0466842
R3980 VSS.n2315 VSS.n31 0.0466842
R3981 VSS.n1611 VSS.n1610 0.0466842
R3982 VSS.n1468 VSS.n484 0.0466842
R3983 VSS.n1307 VSS.n537 0.0466842
R3984 VSS.n1179 VSS.n591 0.0466842
R3985 VSS.n2178 VSS.n2121 0.0466842
R3986 VSS.n1067 VSS.n1066 0.0466842
R3987 VSS VSS.n694 0.0446667
R3988 VSS.n1130 VSS.n606 0.0443158
R3989 VSS.n1258 VSS.n552 0.0443158
R3990 VSS.n1386 VSS.n499 0.0443158
R3991 VSS.n1514 VSS.n431 0.0443158
R3992 VSS.n1553 VSS.n357 0.0443158
R3993 VSS.n2268 VSS.n2267 0.0443158
R3994 VSS.n2104 VSS.n2100 0.0348421
R3995 VSS.n766 VSS 0.0307778
R3996 VSS.n565 VSS 0.0307778
R3997 VSS.n511 VSS 0.0307778
R3998 VSS.n1512 VSS 0.0307778
R3999 VSS.n423 VSS 0.0307778
R4000 VSS.n2242 VSS 0.0307778
R4001 VSS VSS.n2359 0.0307778
R4002 VSS.n2240 VSS 0.0307778
R4003 VSS.n93 VSS.n92 0.0289211
R4004 VSS VSS.n1983 0.0260634
R4005 VSS.n1757 VSS 0.0260634
R4006 VSS.n1685 VSS 0.0260634
R4007 VSS.n311 VSS 0.0260634
R4008 VSS.n923 VSS 0.0260634
R4009 VSS.n958 VSS 0.0260634
R4010 VSS.n2051 VSS.n1983 0.0233169
R4011 VSS.n1757 VSS.n1756 0.0233169
R4012 VSS.n1685 VSS.n1673 0.0233169
R4013 VSS.n888 VSS.n311 0.0233169
R4014 VSS.n924 VSS.n923 0.0233169
R4015 VSS.n959 VSS.n958 0.0233169
R4016 VSS.n2052 VSS.n2051 0.0119085
R4017 VSS.n1756 VSS.n266 0.0119085
R4018 VSS.n1673 VSS.n1671 0.0119085
R4019 VSS.n889 VSS.n888 0.0119085
R4020 VSS.n924 VSS.n831 0.0119085
R4021 VSS.n959 VSS.n767 0.0119085
R4022 VSS.n226 VSS.n54 0.00997368
R4023 VSS.n2047 VSS.n2046 0.00852817
R4024 VSS.n1982 VSS.n1981 0.00852817
R4025 VSS.n1684 VSS.n1682 0.00852817
R4026 VSS.n310 VSS.n285 0.00852817
R4027 VSS.n922 VSS.n877 0.00852817
R4028 VSS.n957 VSS.n814 0.00852817
R4029 VSS.n2149 VSS.n2148 0.00523684
R4030 VSS VSS.n182 0.00383333
R4031 VSS.n2047 VSS 0.0011338
R4032 VSS.n1981 VSS 0.0011338
R4033 VSS VSS.n1684 0.0011338
R4034 VSS VSS.n310 0.0011338
R4035 VSS VSS.n922 0.0011338
R4036 VSS VSS.n957 0.0011338
R4037 OUT.n3 OUT.t3 39.434
R4038 OUT.n0 OUT.t5 39.434
R4039 OUT.n3 OUT.t4 29.3205
R4040 OUT.n0 OUT.t2 29.3205
R4041 OUT.n1 OUT.t1 13.7342
R4042 OUT.n2 OUT.n0 8.09525
R4043 OUT.n1 OUT.t0 6.3271
R4044 OUT OUT.n3 1.09775
R4045 OUT.n3 OUT.n2 1.02275
R4046 OUT.n2 OUT.n1 0.3305
R4047 VCNS.n0 VCNS.t3 40.4718
R4048 VCNS.n2 VCNS.t1 40.4081
R4049 VCNS.n1 VCNS.t2 40.4081
R4050 VCNS.n0 VCNS.t0 40.4081
R4051 VCNS VCNS.n2 1.89975
R4052 VCNS.n1 VCNS.n0 0.06425
R4053 VCNS.n2 VCNS.n1 0.06425
R4054 VCNB.n0 VCNB.t2 40.4718
R4055 VCNB.n2 VCNB.t0 40.4081
R4056 VCNB.n1 VCNB.t3 40.4081
R4057 VCNB.n0 VCNB.t1 40.4081
R4058 VCNB VCNB.n2 1.90056
R4059 VCNB.n1 VCNB.n0 0.06425
R4060 VCNB.n2 VCNB.n1 0.06425
R4061 VCTRL VCTRL.t0 29.2551
C0 a_18489_n1138 OUT 0.058694f
C1 a_11009_2840 VDD 0.454061f
C2 a_14657_n1138 OUT 0.046681f
C3 a_7177_2840 VDD 0.454061f
C4 VDD VCNB 0.115897f
C5 a_18477_2840 VDD 0.298308f
C6 a_3345_2840 VDD 0.454061f
C7 a_14645_2840 VDD 0.298285f
C8 a_n671_n1138 OUT 0.058694f
C9 a_n487_2840 VDD 0.454061f
C10 a_10813_2840 VDD 0.298285f
C11 a_18673_2840 OUT 0.522564f
C12 OUT a_n683_2840 0.198022f
C13 a_6981_2840 VDD 0.298285f
C14 a_n8659_n1230 VCNS 0.1952f
C15 a_7177_2840 a_11009_2840 0.971124f
C16 a_3149_2840 a_3345_2840 0.099479f
C17 a_3149_2840 a_n487_2840 0.072091f
C18 a_14645_2840 a_11009_2840 0.072091f
C19 a_3345_2840 a_7177_2840 0.971124f
C20 a_10813_2840 a_11009_2840 0.099479f
C21 a_10813_2840 a_7177_2840 0.072091f
C22 a_n487_2840 a_3345_2840 0.971124f
C23 a_6981_2840 a_7177_2840 0.099479f
C24 a_18673_2840 VDD 0.282552f
C25 a_6981_2840 a_3345_2840 0.072091f
C26 VDD a_n683_2840 0.298285f
C27 VDD a_n9701_6193 0.406316f
C28 VDD OUT 1.71981f
C29 a_11009_2840 a_14657_n1138 0.058694f
C30 a_11009_2840 a_10825_n1138 0.046681f
C31 a_7177_2840 a_10825_n1138 0.058694f
C32 VDD VCNS 0.199523f
C33 a_7177_2840 a_6993_n1138 0.046681f
C34 a_3345_2840 a_6993_n1138 0.058694f
C35 a_3345_2840 a_3161_n1138 0.046681f
C36 a_n8659_n1230 VCNB 0.205658f
C37 VCTRL a_n9701_6193 0.073173f
C38 a_3149_2840 OUT 0.122036f
C39 a_n487_2840 a_3161_n1138 0.058694f
C40 a_18477_2840 a_18673_2840 0.106065f
C41 a_n487_2840 a_n671_n1138 0.046681f
C42 a_11009_2840 OUT 1.11554f
C43 a_7177_2840 OUT 0.142403f
C44 a_18477_2840 OUT 0.073021f
C45 a_n487_2840 a_n683_2840 0.099479f
C46 a_3345_2840 OUT 0.142403f
C47 a_14645_2840 OUT 0.222712f
C48 a_n487_2840 OUT 1.12692f
C49 a_10813_2840 OUT 0.122036f
C50 a_6981_2840 OUT 0.122036f
C51 a_18673_2840 a_18489_n1138 0.063905f
C52 VDD VCTRL 0.130527f
C53 a_3149_2840 VDD 0.298285f
C54 VCNS VSS 2.63992f
C55 VCNB VSS 2.51968f
C56 OUT VSS 13.7717f
C57 VCTRL VSS 2.27922f
C58 VDD VSS 80.1318f
C59 a_18489_n1138 VSS 0.702283f
C60 a_14657_n1138 VSS 0.709529f
C61 a_10825_n1138 VSS 0.709529f
C62 a_6993_n1138 VSS 0.709529f
C63 a_3161_n1138 VSS 0.709529f
C64 a_n671_n1138 VSS 0.709529f
C65 a_n8659_n1230 VSS 2.37379f
C66 a_18673_2840 VSS 1.21564f
C67 a_11009_2840 VSS 3.67928f
C68 a_7177_2840 VSS 3.67928f
C69 a_18477_2840 VSS 0.393424f
C70 a_3345_2840 VSS 3.67928f
C71 a_14645_2840 VSS 0.393424f
C72 a_n487_2840 VSS 3.6607f
C73 a_10813_2840 VSS 0.393424f
C74 a_6981_2840 VSS 0.393424f
C75 a_3149_2840 VSS 0.393424f
C76 a_n683_2840 VSS 0.393424f
C77 a_n9701_6193 VSS 3.11268f
C78 a_16431_6193 VSS 0.776388f
C79 a_n4208_n141.n0 VSS 0.127578f
C80 a_n4208_n141.n1 VSS 1.58f
C81 a_n4208_n141.n2 VSS 0.69432f
C82 a_n4208_n141.n3 VSS 0.890258f
C83 a_n4208_n141.t4 VSS 0.020224f
C84 a_n4208_n141.t0 VSS 0.052649f
C85 VDD.t14 VSS 0.065802f
C86 VDD.n2 VSS 0.04396f
C87 VDD.t0 VSS 0.09131f
C88 VDD.n3 VSS 0.091175f
C89 VDD.n5 VSS 0.12304f
C90 VDD.t6 VSS 0.065802f
C91 VDD.n8 VSS 0.04396f
C92 VDD.t19 VSS 0.09131f
C93 VDD.n9 VSS 0.091175f
C94 VDD.n11 VSS 0.065116f
C95 VDD.n12 VSS 0.21043f
C96 VDD.t2 VSS 0.065802f
C97 VDD.n15 VSS 0.04396f
C98 VDD.t21 VSS 0.09131f
C99 VDD.n16 VSS 0.091175f
C100 VDD.n18 VSS 0.065116f
C101 VDD.n19 VSS 0.209286f
C102 VDD.t4 VSS 0.065802f
C103 VDD.n22 VSS 0.04396f
C104 VDD.t18 VSS 0.09131f
C105 VDD.n23 VSS 0.091175f
C106 VDD.n25 VSS 0.065116f
C107 VDD.n26 VSS 0.209286f
C108 VDD.t16 VSS 0.065802f
C109 VDD.n29 VSS 0.04396f
C110 VDD.t20 VSS 0.09131f
C111 VDD.n30 VSS 0.091175f
C112 VDD.n32 VSS 0.065116f
C113 VDD.n33 VSS 0.209286f
C114 VDD.t10 VSS 0.065802f
C115 VDD.n36 VSS 0.04396f
C116 VDD.t1 VSS 0.09131f
C117 VDD.n37 VSS 0.091175f
C118 VDD.n39 VSS 0.065116f
C119 VDD.n40 VSS 0.209286f
C120 VDD.t8 VSS 0.065802f
C121 VDD.n41 VSS 0.069914f
C122 VDD.t12 VSS 0.065802f
C123 VDD.n42 VSS 0.073569f
C124 VDD.n43 VSS 0.10713f
C125 VDD.n44 VSS 0.268705f
C126 a_n8471_219.n0 VSS 2.95013f
C127 a_n8471_219.n1 VSS 1.11094f
C128 a_n8471_219.n2 VSS 1.43208f
C129 a_n8471_219.n3 VSS 0.328251f
C130 a_n8471_219.t3 VSS 0.036811f
C131 a_n8471_219.t0 VSS 0.038078f
C132 a_n8471_219.t2 VSS 0.012483f
C133 a_n8471_219.t8 VSS 0.012265f
C134 a_n8471_219.t6 VSS 0.029697f
C135 a_n8471_219.t9 VSS 0.010598f
C136 a_n8471_219.t11 VSS 0.010598f
C137 a_n8471_219.t10 VSS 0.010598f
C138 a_n8471_219.t5 VSS 0.010598f
C139 a_n8471_219.t7 VSS 0.010598f
C140 a_n8471_219.t4 VSS 0.022976f
C141 a_n8471_219.n4 VSS 0.365741f
.ends

