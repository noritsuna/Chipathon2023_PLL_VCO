* Extracted by KLayout with GF180MCU LVS runset on : 08/01/2024 22:35

.SUBCKT TOP VSS VCNS VCNB vctrl OUT
R$2 VSS \$33 VSS 227500 ppolyf_u L=520U W=0.8U
M$5 VSS VCNS \$12 VSS nfet_03v3_dn L=0.33U W=8U AS=2.78P AD=2.78P PS=12.78U
+ PD=12.78U
M$9 \$13 VCNB \$12 VSS nfet_03v3_dn L=0.33U W=8U AS=2.78P AD=2.78P PS=12.78U
+ PD=12.78U
M$13 \$33 vctrl \$13 VSS nfet_03v3_dn L=0.33U W=0.8U AS=0.488P AD=0.488P
+ PS=2.82U PD=2.82U
M$14 \$1 \$13 \$6 \$1 pfet_03v3 L=0.33U W=1.8U AS=1.17P AD=1.17P PS=4.9U PD=4.9U
M$15 \$32 OUT \$I159 \$1 pfet_03v3 L=0.33U W=3.6U AS=2.34P AD=2.34P PS=8.5U
+ PD=8.5U
M$16 \$I55 \$I63 \$I171 \$1 pfet_03v3 L=0.33U W=3.6U AS=2.34P AD=2.34P PS=8.5U
+ PD=8.5U
M$17 \$I63 OUT \$I183 \$1 pfet_03v3 L=0.33U W=3.6U AS=2.34P AD=2.34P PS=8.5U
+ PD=8.5U
M$18 \$I56 \$I55 \$I195 \$1 pfet_03v3 L=0.33U W=3.6U AS=2.34P AD=2.34P PS=8.5U
+ PD=8.5U
M$19 \$I57 \$I56 \$I207 \$1 pfet_03v3 L=0.33U W=3.6U AS=2.34P AD=2.34P PS=8.5U
+ PD=8.5U
M$20 OUT \$I57 \$I219 \$1 pfet_03v3 L=0.33U W=3.6U AS=2.34P AD=2.34P PS=8.5U
+ PD=8.5U
M$21 \$1 \$13 \$13 \$1 pfet_03v3 L=0.33U W=1.8U AS=1.17P AD=1.17P PS=4.9U
+ PD=4.9U
M$22 \$1 \$13 \$I159 \$1 pfet_03v3 L=0.33U W=1.8U AS=1.17P AD=1.17P PS=4.9U
+ PD=4.9U
M$23 \$1 \$13 \$I171 \$1 pfet_03v3 L=0.33U W=1.8U AS=1.17P AD=1.17P PS=4.9U
+ PD=4.9U
M$24 \$1 \$13 \$I183 \$1 pfet_03v3 L=0.33U W=1.8U AS=1.17P AD=1.17P PS=4.9U
+ PD=4.9U
M$25 \$1 \$13 \$I195 \$1 pfet_03v3 L=0.33U W=1.8U AS=1.17P AD=1.17P PS=4.9U
+ PD=4.9U
M$26 \$1 \$13 \$I207 \$1 pfet_03v3 L=0.33U W=1.8U AS=1.17P AD=1.17P PS=4.9U
+ PD=4.9U
M$27 \$1 \$13 \$I219 \$1 pfet_03v3 L=0.33U W=1.8U AS=1.17P AD=1.17P PS=4.9U
+ PD=4.9U
M$28 VSS \$6 \$6 VSS nfet_03v3_dn L=0.33U W=0.7U AS=0.427P AD=0.427P PS=2.62U
+ PD=2.62U
M$29 VSS \$6 \$I155 VSS nfet_03v3_dn L=0.33U W=0.7U AS=0.427P AD=0.427P
+ PS=2.62U PD=2.62U
M$30 VSS \$6 \$I167 VSS nfet_03v3_dn L=0.33U W=0.7U AS=0.427P AD=0.427P
+ PS=2.62U PD=2.62U
M$31 VSS \$6 \$I179 VSS nfet_03v3_dn L=0.33U W=0.7U AS=0.427P AD=0.427P
+ PS=2.62U PD=2.62U
M$32 VSS \$6 \$I191 VSS nfet_03v3_dn L=0.33U W=0.7U AS=0.427P AD=0.427P
+ PS=2.62U PD=2.62U
M$33 VSS \$6 \$I203 VSS nfet_03v3_dn L=0.33U W=0.7U AS=0.427P AD=0.427P
+ PS=2.62U PD=2.62U
M$34 VSS \$6 \$I215 VSS nfet_03v3_dn L=0.33U W=0.7U AS=0.427P AD=0.427P
+ PS=2.62U PD=2.62U
M$35 \$32 OUT \$I155 VSS nfet_03v3_dn L=0.33U W=1.4U AS=0.854P AD=0.854P
+ PS=4.02U PD=4.02U
M$36 \$I55 \$I63 \$I167 VSS nfet_03v3_dn L=0.33U W=1.4U AS=0.854P AD=0.854P
+ PS=4.02U PD=4.02U
M$37 \$I63 OUT \$I179 VSS nfet_03v3_dn L=0.33U W=1.4U AS=0.854P AD=0.854P
+ PS=4.02U PD=4.02U
M$38 \$I56 \$I55 \$I191 VSS nfet_03v3_dn L=0.33U W=1.4U AS=0.854P AD=0.854P
+ PS=4.02U PD=4.02U
M$39 \$I57 \$I56 \$I203 VSS nfet_03v3_dn L=0.33U W=1.4U AS=0.854P AD=0.854P
+ PS=4.02U PD=4.02U
M$40 OUT \$I57 \$I215 VSS nfet_03v3_dn L=0.33U W=1.4U AS=0.854P AD=0.854P
+ PS=4.02U PD=4.02U
.ENDS TOP
