* NGSPICE file created from TOP.ext - technology: gf180mcuD

.subckt TOP VDD VCTRL OUT VCNB VCNS VSS
X0 VDD.t20 a_n8471_219.t5 a_3149_2840 VDD.t19 pfet_03v3 ad=0.585p pd=3.1u as=0.585p ps=3.1u w=0.9u l=0.33u
X1 VSS.t29 a_n4208_n141.t3 a_n671_n1138 VSS.t28 nfet_03v3 ad=0.2646p pd=2.1u as=0.2646p ps=2.1u w=0.42u l=0.33u
X2 OUT.t0 a_11009_2840 a_14657_n1138 VSS.t5 nfet_03v3 ad=0.5124p pd=2.9u as=0.5124p ps=2.9u w=0.84u l=0.33u
X3 a_7177_2840 a_3345_2840 a_6981_2840 VDD.t4 pfet_03v3 ad=1.17p pd=4.9u as=1.17p ps=4.9u w=1.8u l=0.33u
X4 VSS.t10 VCNS.t0 a_n8659_n1230 VSS.t9 nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.33u
X5 VSS.t34 a_16431_6193 VSS.t30 ppolyf_u r_width=0.8u r_length=0.13m
X6 a_n8471_219.t1 VCNB.t0 a_n8659_n1230 VSS.t4 nfet_03v3 ad=0.52p pd=2.52u as=1.22p ps=5.22u w=2u l=0.33u
X7 VDD.t18 a_n8471_219.t6 a_18477_2840 VDD.t17 pfet_03v3 ad=0.585p pd=3.1u as=0.585p ps=3.1u w=0.9u l=0.33u
X8 VSS.t15 VCNS.t1 a_n8659_n1230 VSS.t14 nfet_03v3 ad=0.52p pd=2.52u as=1.22p ps=5.22u w=2u l=0.33u
X9 VDD.t16 a_n8471_219.t3 a_n8471_219.t4 VDD.t15 pfet_03v3 ad=0.585p pd=3.1u as=0.585p ps=3.1u w=0.9u l=0.33u
X10 VDD.t14 a_n8471_219.t7 a_n683_2840 VDD.t13 pfet_03v3 ad=0.585p pd=3.1u as=0.585p ps=3.1u w=0.9u l=0.33u
X11 a_11009_2840 a_7177_2840 a_10813_2840 VDD.t3 pfet_03v3 ad=1.17p pd=4.9u as=1.17p ps=4.9u w=1.8u l=0.33u
X12 a_3345_2840 a_n487_2840 a_3149_2840 VDD.t2 pfet_03v3 ad=1.17p pd=4.9u as=1.17p ps=4.9u w=1.8u l=0.33u
X13 a_n4208_n141.t2 a_n8471_219.t8 VDD.t12 VDD.t11 pfet_03v3 ad=0.585p pd=3.1u as=0.585p ps=3.1u w=0.9u l=0.33u
X14 a_n487_2840 OUT.t2 a_n671_n1138 VSS.t1 nfet_03v3 ad=0.5124p pd=2.9u as=0.5124p ps=2.9u w=0.84u l=0.33u
X15 a_7177_2840 a_3345_2840 a_6993_n1138 VSS.t33 nfet_03v3 ad=0.5124p pd=2.9u as=0.5124p ps=2.9u w=0.84u l=0.33u
X16 a_n8471_219.t0 VCTRL.t0 a_n9701_6193 VSS.t0 nfet_03v3 ad=0.488p pd=2.82u as=0.488p ps=2.82u w=0.8u l=0.33u
X17 a_18673_2840 OUT.t3 a_18477_2840 VDD.t21 pfet_03v3 ad=1.17p pd=4.9u as=1.17p ps=4.9u w=1.8u l=0.33u
X18 a_18673_2840 OUT.t4 a_18489_n1138 VSS.t13 nfet_03v3 ad=0.5124p pd=2.9u as=0.5124p ps=2.9u w=0.84u l=0.33u
X19 VSS.t27 a_n4208_n141.t4 a_18489_n1138 VSS.t26 nfet_03v3 ad=0.2646p pd=2.1u as=0.2646p ps=2.1u w=0.42u l=0.33u
X20 a_n487_2840 OUT.t5 a_n683_2840 VDD.t1 pfet_03v3 ad=1.17p pd=4.9u as=1.17p ps=4.9u w=1.8u l=0.33u
X21 a_n8659_n1230 VCNS.t2 VSS.t3 VSS.t2 nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.33u
X22 VDD.t10 a_n8471_219.t9 a_14645_2840 VDD.t9 pfet_03v3 ad=0.585p pd=3.1u as=0.585p ps=3.1u w=0.9u l=0.33u
X23 VSS.t25 a_n4208_n141.t5 a_14657_n1138 VSS.t24 nfet_03v3 ad=0.2646p pd=2.1u as=0.2646p ps=2.1u w=0.42u l=0.33u
X24 VSS.t23 a_n4208_n141.t6 a_3161_n1138 VSS.t22 nfet_03v3 ad=0.2646p pd=2.1u as=0.2646p ps=2.1u w=0.42u l=0.33u
X25 VDD.t8 a_n8471_219.t10 a_6981_2840 VDD.t7 pfet_03v3 ad=0.585p pd=3.1u as=0.585p ps=3.1u w=0.9u l=0.33u
X26 a_n8471_219.t2 VCNB.t1 a_n8659_n1230 VSS.t8 nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.33u
X27 a_n4208_n141.t1 a_n4208_n141.t0 VSS.t21 VSS.t20 nfet_03v3 ad=0.2646p pd=2.1u as=0.2646p ps=2.1u w=0.42u l=0.33u
X28 a_11009_2840 a_7177_2840 a_10825_n1138 VSS.t32 nfet_03v3 ad=0.5124p pd=2.9u as=0.5124p ps=2.9u w=0.84u l=0.33u
X29 VSS.t19 a_n4208_n141.t7 a_6993_n1138 VSS.t18 nfet_03v3 ad=0.2646p pd=2.1u as=0.2646p ps=2.1u w=0.42u l=0.33u
X30 a_n8659_n1230 VCNB.t2 a_n8471_219.t2 VSS.t11 nfet_03v3 ad=1.22p pd=5.22u as=0.52p ps=2.52u w=2u l=0.33u
X31 a_n8659_n1230 VCNS.t3 VSS.t7 VSS.t6 nfet_03v3 ad=1.22p pd=5.22u as=0.52p ps=2.52u w=2u l=0.33u
X32 a_3345_2840 a_n487_2840 a_3161_n1138 VSS.t31 nfet_03v3 ad=0.5124p pd=2.9u as=0.5124p ps=2.9u w=0.84u l=0.33u
X33 VSS.t17 a_n4208_n141.t8 a_10825_n1138 VSS.t16 nfet_03v3 ad=0.2646p pd=2.1u as=0.2646p ps=2.1u w=0.42u l=0.33u
X34 a_n9701_6193 a_16431_6193 VSS.t30 ppolyf_u r_width=0.8u r_length=0.13m
X35 VDD.t6 a_n8471_219.t11 a_10813_2840 VDD.t5 pfet_03v3 ad=0.585p pd=3.1u as=0.585p ps=3.1u w=0.9u l=0.33u
X36 a_n8659_n1230 VCNB.t3 a_n8471_219.t1 VSS.t12 nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.33u
X37 OUT.t1 a_11009_2840 a_14645_2840 VDD.t0 pfet_03v3 ad=1.17p pd=4.9u as=1.17p ps=4.9u w=1.8u l=0.33u
R0 a_n8471_219.n1 a_n8471_219.t6 31.1854
R1 a_n8471_219.n0 a_n8471_219.t8 30.4809
R2 a_n8471_219.n0 a_n8471_219.t7 29.7468
R3 a_n8471_219.n0 a_n8471_219.t5 29.7468
R4 a_n8471_219.n2 a_n8471_219.t10 29.7468
R5 a_n8471_219.n2 a_n8471_219.t11 29.7468
R6 a_n8471_219.n1 a_n8471_219.t9 29.7468
R7 a_n8471_219.n3 a_n8471_219.t3 28.2414
R8 a_n8471_219.n0 a_n8471_219.t0 11.7439
R9 a_n8471_219.n3 a_n8471_219.t4 8.52921
R10 a_n8471_219.t1 a_n8471_219.n4 4.56638
R11 a_n8471_219.n4 a_n8471_219.t2 4.38259
R12 a_n8471_219.n4 a_n8471_219.n0 3.5234
R13 a_n8471_219.n0 a_n8471_219.n2 2.8778
R14 a_n8471_219.n2 a_n8471_219.n1 2.8778
R15 a_n8471_219.n0 a_n8471_219.n3 2.4541
R16 VDD.n2 VDD.t17 589.355
R17 VDD.n8 VDD.t9 589.355
R18 VDD.n15 VDD.t5 589.355
R19 VDD.n22 VDD.t7 589.355
R20 VDD.n29 VDD.t19 589.355
R21 VDD.n36 VDD.t13 589.355
R22 VDD.n42 VDD.t15 589.355
R23 VDD.n41 VDD.t11 589.355
R24 VDD.n3 VDD.t21 419.211
R25 VDD.n9 VDD.t0 419.211
R26 VDD.n16 VDD.t3 419.211
R27 VDD.n23 VDD.t4 419.211
R28 VDD.n30 VDD.t2 419.211
R29 VDD.n37 VDD.t1 419.211
R30 VDD.n42 VDD.t16 8.52192
R31 VDD.n41 VDD.t12 8.52192
R32 VDD.n2 VDD.t18 8.46717
R33 VDD.n8 VDD.t10 8.46717
R34 VDD.n15 VDD.t6 8.46717
R35 VDD.n22 VDD.t8 8.46717
R36 VDD.n29 VDD.t20 8.46717
R37 VDD.n36 VDD.t14 8.46717
R38 VDD.n4 VDD.n1 4.5005
R39 VDD.n1 VDD.n0 4.5005
R40 VDD.n4 VDD.n3 4.5005
R41 VDD.n3 VDD.n0 4.5005
R42 VDD.n10 VDD.n7 4.5005
R43 VDD.n7 VDD.n6 4.5005
R44 VDD.n10 VDD.n9 4.5005
R45 VDD.n9 VDD.n6 4.5005
R46 VDD.n17 VDD.n14 4.5005
R47 VDD.n14 VDD.n13 4.5005
R48 VDD.n17 VDD.n16 4.5005
R49 VDD.n16 VDD.n13 4.5005
R50 VDD.n24 VDD.n21 4.5005
R51 VDD.n21 VDD.n20 4.5005
R52 VDD.n24 VDD.n23 4.5005
R53 VDD.n23 VDD.n20 4.5005
R54 VDD.n31 VDD.n28 4.5005
R55 VDD.n28 VDD.n27 4.5005
R56 VDD.n31 VDD.n30 4.5005
R57 VDD.n30 VDD.n27 4.5005
R58 VDD.n38 VDD.n35 4.5005
R59 VDD.n35 VDD.n34 4.5005
R60 VDD.n38 VDD.n37 4.5005
R61 VDD.n37 VDD.n34 4.5005
R62 VDD.n44 VDD.n43 4.06871
R63 VDD VDD.n5 3.40475
R64 VDD.n12 VDD.n11 2.70462
R65 VDD.n19 VDD.n18 2.70462
R66 VDD.n26 VDD.n25 2.70462
R67 VDD.n33 VDD.n32 2.70462
R68 VDD.n40 VDD.n39 2.70462
R69 VDD VDD.n44 0.777875
R70 VDD.n12 VDD 0.737375
R71 VDD.n19 VDD 0.7265
R72 VDD.n26 VDD 0.7265
R73 VDD.n33 VDD 0.7265
R74 VDD.n40 VDD 0.7265
R75 VDD.n44 VDD 0.7265
R76 VDD VDD.n12 0.7115
R77 VDD VDD.n19 0.7115
R78 VDD VDD.n26 0.7115
R79 VDD VDD.n33 0.7115
R80 VDD VDD.n40 0.7115
R81 VDD.n43 VDD.n42 0.181952
R82 VDD.n43 VDD.n41 0.146702
R83 VDD.n5 VDD.n4 0.024117
R84 VDD.n11 VDD.n10 0.024117
R85 VDD.n18 VDD.n17 0.024117
R86 VDD.n25 VDD.n24 0.024117
R87 VDD.n32 VDD.n31 0.024117
R88 VDD.n39 VDD.n38 0.024117
R89 VDD.n5 VDD.n0 0.0237979
R90 VDD.n11 VDD.n6 0.0237979
R91 VDD.n18 VDD.n13 0.0237979
R92 VDD.n25 VDD.n20 0.0237979
R93 VDD.n32 VDD.n27 0.0237979
R94 VDD.n39 VDD.n34 0.0237979
R95 VDD.n2 VDD.n1 0.020375
R96 VDD.n3 VDD.n2 0.020375
R97 VDD.n8 VDD.n7 0.020375
R98 VDD.n9 VDD.n8 0.020375
R99 VDD.n15 VDD.n14 0.020375
R100 VDD.n16 VDD.n15 0.020375
R101 VDD.n22 VDD.n21 0.020375
R102 VDD.n23 VDD.n22 0.020375
R103 VDD.n29 VDD.n28 0.020375
R104 VDD.n30 VDD.n29 0.020375
R105 VDD.n36 VDD.n35 0.020375
R106 VDD.n37 VDD.n36 0.020375
R107 a_n4208_n141.n2 a_n4208_n141.t4 26.5147
R108 a_n4208_n141.n1 a_n4208_n141.t3 25.076
R109 a_n4208_n141.n1 a_n4208_n141.t6 25.076
R110 a_n4208_n141.n3 a_n4208_n141.t7 25.076
R111 a_n4208_n141.n3 a_n4208_n141.t8 25.076
R112 a_n4208_n141.n2 a_n4208_n141.t5 25.076
R113 a_n4208_n141.n0 a_n4208_n141.t0 23.009
R114 a_n4208_n141.n0 a_n4208_n141.t1 12.3005
R115 a_n4208_n141.t2 a_n4208_n141.n1 11.2556
R116 a_n4208_n141.n1 a_n4208_n141.n0 3.08843
R117 a_n4208_n141.n1 a_n4208_n141.n3 2.8778
R118 a_n4208_n141.n3 a_n4208_n141.n2 2.8778
R119 VSS.n2271 VSS.n2231 168832
R120 VSS.n1479 VSS.n188 136590
R121 VSS.n741 VSS.n740 134875
R122 VSS.n1485 VSS.n1484 134875
R123 VSS.n1483 VSS.n1482 134875
R124 VSS.n1481 VSS.n1480 134875
R125 VSS.n741 VSS.n513 126750
R126 VSS.n1484 VSS.n1483 126750
R127 VSS.n1482 VSS.n1481 126750
R128 VSS.n1480 VSS.n1479 126750
R129 VSS.n1913 VSS.n188 65268.1
R130 VSS.n2271 VSS.n2270 63487.1
R131 VSS.n2028 VSS.n2027 23007.5
R132 VSS.n224 VSS.n223 17472.4
R133 VSS.n1790 VSS.n222 13029.1
R134 VSS.n2231 VSS.n2230 11767.2
R135 VSS.n2230 VSS.n80 11262.4
R136 VSS.n2056 VSS.n2055 6332.65
R137 VSS.n2027 VSS.n130 5968.01
R138 VSS.n1991 VSS.n130 5872.22
R139 VSS.n2270 VSS.n2232 5104.34
R140 VSS.n222 VSS.n117 4375.37
R141 VSS.n744 VSS.n741 3636.7
R142 VSS.n1484 VSS.n117 3636.7
R143 VSS.n1482 VSS.n117 3636.7
R144 VSS.n1480 VSS.n117 3636.7
R145 VSS.n1682 VSS.n1655 2950.24
R146 VSS.n1682 VSS.n224 2950.24
R147 VSS.n1655 VSS.n267 2950.24
R148 VSS.n849 VSS.n267 2950.24
R149 VSS.n849 VSS.n117 2950.24
R150 VSS.n744 VSS.n518 2950.24
R151 VSS.n1790 VSS.n224 2338.06
R152 VSS.n1707 VSS.n117 1959.56
R153 VSS.n1024 VSS.n117 1959.56
R154 VSS.n1059 VSS.n117 1959.56
R155 VSS.n1094 VSS.n117 1959.56
R156 VSS.n1129 VSS.n117 1959.56
R157 VSS.n188 VSS.n117 1872.67
R158 VSS.n1996 VSS.t20 1362.36
R159 VSS.t30 VSS.n2057 1272.15
R160 VSS.n2367 VSS.t0 1191.42
R161 VSS.n456 VSS.t24 948.962
R162 VSS.n376 VSS.t18 948.962
R163 VSS.n153 VSS.t28 948.962
R164 VSS.n375 VSS.t22 948.962
R165 VSS.n379 VSS.t16 948.962
R166 VSS.n666 VSS.t26 948.962
R167 VSS.n456 VSS.t5 873.535
R168 VSS.n376 VSS.t33 873.535
R169 VSS.n153 VSS.t1 873.535
R170 VSS.n375 VSS.t31 873.535
R171 VSS.n379 VSS.t32 873.535
R172 VSS.n666 VSS.t13 873.535
R173 VSS.n223 VSS.n117 814.926
R174 VSS.n2331 VSS.t4 782.77
R175 VSS.n550 VSS.n545 781.367
R176 VSS.n2316 VSS.t14 769.106
R177 VSS.n2269 VSS.n2233 583.484
R178 VSS.n2263 VSS.n2233 583.484
R179 VSS.n2263 VSS.n2262 583.484
R180 VSS.n2262 VSS.n2261 583.484
R181 VSS.n2261 VSS.n2244 583.484
R182 VSS.n2255 VSS.n2244 583.484
R183 VSS.n2255 VSS.n2254 583.484
R184 VSS.n2254 VSS.n49 583.484
R185 VSS.n1432 VSS.n1409 534.539
R186 VSS.n1432 VSS.n1431 534.539
R187 VSS.n1431 VSS.n1430 534.539
R188 VSS.n1430 VSS.n1410 534.539
R189 VSS.n1424 VSS.n1410 534.539
R190 VSS.n1424 VSS.n1423 534.539
R191 VSS.n1301 VSS.n1255 534.539
R192 VSS.n1301 VSS.n1300 534.539
R193 VSS.n1300 VSS.n1299 534.539
R194 VSS.n1299 VSS.n1278 534.539
R195 VSS.n1293 VSS.n1278 534.539
R196 VSS.n1293 VSS.n1292 534.539
R197 VSS.n1388 VSS.n1250 534.539
R198 VSS.n1388 VSS.n1387 534.539
R199 VSS.n1387 VSS.n1386 534.539
R200 VSS.n1386 VSS.n1251 534.539
R201 VSS.n1380 VSS.n1251 534.539
R202 VSS.n1380 VSS.n1379 534.539
R203 VSS.n1219 VSS.n1218 534.539
R204 VSS.n1220 VSS.n1219 534.539
R205 VSS.n1220 VSS.n453 534.539
R206 VSS.n1227 VSS.n453 534.539
R207 VSS.n1228 VSS.n1227 534.539
R208 VSS.n1229 VSS.n1228 534.539
R209 VSS.n693 VSS.n670 534.539
R210 VSS.n693 VSS.n692 534.539
R211 VSS.n692 VSS.n691 534.539
R212 VSS.n691 VSS.n671 534.539
R213 VSS.n685 VSS.n671 534.539
R214 VSS.n685 VSS.n684 534.539
R215 VSS.n1965 VSS.n1964 534.539
R216 VSS.n1966 VSS.n1965 534.539
R217 VSS.n1966 VSS.n150 534.539
R218 VSS.n1973 VSS.n150 534.539
R219 VSS.n1974 VSS.n1973 534.539
R220 VSS.n1975 VSS.n1974 534.539
R221 VSS.t8 VSS.t11 519.268
R222 VSS.t12 VSS.t8 519.268
R223 VSS.t4 VSS.t12 519.268
R224 VSS.n2302 VSS.n49 513.466
R225 VSS.t9 VSS.t6 510.158
R226 VSS.t2 VSS.t9 510.158
R227 VSS.t14 VSS.t2 510.158
R228 VSS.n833 VSS.n117 475.276
R229 VSS.n901 VSS.n117 475.276
R230 VSS.n968 VSS.n117 475.276
R231 VSS.n1699 VSS.n117 475.276
R232 VSS.n2058 VSS.t30 461.793
R233 VSS.n2336 VSS.n28 456.781
R234 VSS.n2336 VSS.n2335 456.781
R235 VSS.n2335 VSS.n2334 456.781
R236 VSS.n2334 VSS.n33 456.781
R237 VSS.n2328 VSS.n33 456.781
R238 VSS.n2328 VSS.n2327 456.781
R239 VSS.n2327 VSS.n2326 456.781
R240 VSS.n2326 VSS.n37 456.781
R241 VSS.n2320 VSS.n37 456.781
R242 VSS.n2320 VSS.n2319 456.781
R243 VSS.n2319 VSS.n2318 456.781
R244 VSS.n2318 VSS.n41 456.781
R245 VSS.n2312 VSS.n41 456.781
R246 VSS.n2312 VSS.n2311 456.781
R247 VSS.n2311 VSS.n2310 456.781
R248 VSS.n2310 VSS.n45 456.781
R249 VSS.n2304 VSS.n45 456.781
R250 VSS.n2304 VSS.n2303 456.781
R251 VSS.n2270 VSS.n2269 425.943
R252 VSS.n744 VSS.n521 364.974
R253 VSS.n1493 VSS.n117 364.974
R254 VSS.n1531 VSS.n117 364.974
R255 VSS.n1569 VSS.n117 364.974
R256 VSS.n1595 VSS.n117 364.974
R257 VSS.n1888 VSS.n117 364.974
R258 VSS.n2224 VSS.n80 354.031
R259 VSS.n2224 VSS.n2223 354.031
R260 VSS.n2223 VSS.n2222 354.031
R261 VSS.n2222 VSS.n2201 354.031
R262 VSS.n2216 VSS.n2201 354.031
R263 VSS.n2057 VSS.n2056 350.44
R264 VSS.n2216 VSS.n20 341.639
R265 VSS.n2342 VSS.n28 326.632
R266 VSS.n2372 VSS.n2371 325.978
R267 VSS.n2371 VSS.n2370 325.978
R268 VSS.n2370 VSS.n11 325.978
R269 VSS.n2363 VSS.n11 325.978
R270 VSS.n2363 VSS.n2362 325.978
R271 VSS.n2362 VSS.n2361 325.978
R272 VSS.n2361 VSS.n16 325.978
R273 VSS.n2355 VSS.n16 325.978
R274 VSS.n2355 VSS.n2354 325.978
R275 VSS.n2354 VSS.n2353 325.978
R276 VSS.n2344 VSS.n2343 325.978
R277 VSS.n2343 VSS.n2342 325.978
R278 VSS.n1775 VSS.n229 316.457
R279 VSS.n1781 VSS.n229 316.457
R280 VSS.n1782 VSS.n1781 316.457
R281 VSS.n1783 VSS.n1782 316.457
R282 VSS.n1783 VSS.n225 316.457
R283 VSS.n1789 VSS.n225 316.457
R284 VSS.n1792 VSS.n1791 316.457
R285 VSS.n1792 VSS.n218 316.457
R286 VSS.n1798 VSS.n218 316.457
R287 VSS.n1799 VSS.n1798 316.457
R288 VSS.n1800 VSS.n1799 316.457
R289 VSS.n1800 VSS.n214 316.457
R290 VSS.n1806 VSS.n214 316.457
R291 VSS.n1807 VSS.n1806 316.457
R292 VSS.n1808 VSS.n1807 316.457
R293 VSS.n1853 VSS.n1852 316.457
R294 VSS.n1852 VSS.n1851 316.457
R295 VSS.n1851 VSS.n1813 316.457
R296 VSS.n1845 VSS.n1813 316.457
R297 VSS.n1845 VSS.n1844 316.457
R298 VSS.n1844 VSS.n1843 316.457
R299 VSS.n1843 VSS.n1817 316.457
R300 VSS.n1837 VSS.n1817 316.457
R301 VSS.n1837 VSS.n1836 316.457
R302 VSS.n1836 VSS.n1835 316.457
R303 VSS.n1835 VSS.n1821 316.457
R304 VSS.n1829 VSS.n1821 316.457
R305 VSS.n1829 VSS.n1828 316.457
R306 VSS.n1828 VSS.n1827 316.457
R307 VSS.n1827 VSS.n131 316.457
R308 VSS.n2026 VSS.n132 316.457
R309 VSS.n2020 VSS.n132 316.457
R310 VSS.n2020 VSS.n2019 316.457
R311 VSS.n2019 VSS.n2018 316.457
R312 VSS.n2137 VSS.n98 310.856
R313 VSS.n1423 VSS.n156 307.361
R314 VSS.n1292 VSS.n358 307.361
R315 VSS.n1379 VSS.n1378 307.361
R316 VSS.n1229 VSS.n447 307.361
R317 VSS.n684 VSS.n458 307.361
R318 VSS.n1975 VSS.n138 307.361
R319 VSS.n1409 VSS.n358 304.688
R320 VSS.n1378 VSS.n1255 304.688
R321 VSS.n1250 VSS.n447 304.688
R322 VSS.n1218 VSS.n458 304.688
R323 VSS.n670 VSS.n654 304.688
R324 VSS.n1964 VSS.n156 304.688
R325 VSS.n2002 VSS.n2001 302.748
R326 VSS.n2001 VSS.n2000 302.748
R327 VSS.n2000 VSS.n1993 302.748
R328 VSS.n1993 VSS.n70 302.748
R329 VSS.n2283 VSS.n70 302.748
R330 VSS.n2283 VSS.n2282 302.748
R331 VSS.n2118 VSS.n98 301.029
R332 VSS.n2018 VSS.n138 287.976
R333 VSS.n733 VSS.n522 278.851
R334 VSS.n733 VSS.n732 278.851
R335 VSS.n732 VSS.n731 278.851
R336 VSS.n731 VSS.n638 278.851
R337 VSS.n725 VSS.n638 278.851
R338 VSS.n725 VSS.n724 278.851
R339 VSS.n724 VSS.n723 278.851
R340 VSS.n723 VSS.n642 278.851
R341 VSS.n717 VSS.n642 278.851
R342 VSS.n717 VSS.n716 278.851
R343 VSS.n716 VSS.n715 278.851
R344 VSS.n715 VSS.n646 278.851
R345 VSS.n709 VSS.n646 278.851
R346 VSS.n709 VSS.n708 278.851
R347 VSS.n708 VSS.n707 278.851
R348 VSS.n707 VSS.n650 278.851
R349 VSS.n550 VSS.n517 278.373
R350 VSS.n745 VSS.n517 278.373
R351 VSS.n2184 VSS.n2140 277.659
R352 VSS.n2178 VSS.n2140 277.659
R353 VSS.n2178 VSS.n2177 277.659
R354 VSS.n2177 VSS.n2176 277.659
R355 VSS.n2176 VSS.n2163 277.659
R356 VSS.n2165 VSS.n2163 277.659
R357 VSS.n2165 VSS.n78 277.659
R358 VSS.n2273 VSS.n2272 277.659
R359 VSS.n2273 VSS.n71 277.659
R360 VSS.n2280 VSS.n72 277.659
R361 VSS.n72 VSS.n60 277.659
R362 VSS.n1472 VSS.n330 270.495
R363 VSS.n1472 VSS.n1471 270.495
R364 VSS.n1471 VSS.n1470 270.495
R365 VSS.n1470 VSS.n342 270.495
R366 VSS.n1464 VSS.n342 270.495
R367 VSS.n1464 VSS.n1463 270.495
R368 VSS.n1463 VSS.n1462 270.495
R369 VSS.n1462 VSS.n346 270.495
R370 VSS.n1456 VSS.n346 270.495
R371 VSS.n1456 VSS.n1455 270.495
R372 VSS.n1455 VSS.n1454 270.495
R373 VSS.n1454 VSS.n350 270.495
R374 VSS.n1448 VSS.n350 270.495
R375 VSS.n1448 VSS.n1447 270.495
R376 VSS.n1447 VSS.n1446 270.495
R377 VSS.n1446 VSS.n354 270.495
R378 VSS.n1345 VSS.n328 270.495
R379 VSS.n1346 VSS.n1345 270.495
R380 VSS.n1347 VSS.n1346 270.495
R381 VSS.n1347 VSS.n1327 270.495
R382 VSS.n1353 VSS.n1327 270.495
R383 VSS.n1354 VSS.n1353 270.495
R384 VSS.n1355 VSS.n1354 270.495
R385 VSS.n1355 VSS.n1323 270.495
R386 VSS.n1361 VSS.n1323 270.495
R387 VSS.n1362 VSS.n1361 270.495
R388 VSS.n1363 VSS.n1362 270.495
R389 VSS.n1363 VSS.n1319 270.495
R390 VSS.n1369 VSS.n1319 270.495
R391 VSS.n1370 VSS.n1369 270.495
R392 VSS.n1371 VSS.n1370 270.495
R393 VSS.n1371 VSS.n1256 270.495
R394 VSS.n414 VSS.n326 270.495
R395 VSS.n414 VSS.n400 270.495
R396 VSS.n420 VSS.n400 270.495
R397 VSS.n421 VSS.n420 270.495
R398 VSS.n422 VSS.n421 270.495
R399 VSS.n422 VSS.n396 270.495
R400 VSS.n428 VSS.n396 270.495
R401 VSS.n429 VSS.n428 270.495
R402 VSS.n430 VSS.n429 270.495
R403 VSS.n430 VSS.n392 270.495
R404 VSS.n436 VSS.n392 270.495
R405 VSS.n437 VSS.n436 270.495
R406 VSS.n438 VSS.n437 270.495
R407 VSS.n438 VSS.n388 270.495
R408 VSS.n445 VSS.n388 270.495
R409 VSS.n446 VSS.n445 270.495
R410 VSS.n1168 VSS.n486 270.495
R411 VSS.n1174 VSS.n486 270.495
R412 VSS.n1175 VSS.n1174 270.495
R413 VSS.n1176 VSS.n1175 270.495
R414 VSS.n1176 VSS.n482 270.495
R415 VSS.n1182 VSS.n482 270.495
R416 VSS.n1183 VSS.n1182 270.495
R417 VSS.n1184 VSS.n1183 270.495
R418 VSS.n1184 VSS.n478 270.495
R419 VSS.n1190 VSS.n478 270.495
R420 VSS.n1191 VSS.n1190 270.495
R421 VSS.n1192 VSS.n1191 270.495
R422 VSS.n1192 VSS.n474 270.495
R423 VSS.n1199 VSS.n474 270.495
R424 VSS.n1200 VSS.n1199 270.495
R425 VSS.n1201 VSS.n1200 270.495
R426 VSS.n1914 VSS.n184 270.495
R427 VSS.n1920 VSS.n184 270.495
R428 VSS.n1921 VSS.n1920 270.495
R429 VSS.n1922 VSS.n1921 270.495
R430 VSS.n1922 VSS.n180 270.495
R431 VSS.n1928 VSS.n180 270.495
R432 VSS.n1929 VSS.n1928 270.495
R433 VSS.n1930 VSS.n1929 270.495
R434 VSS.n1930 VSS.n176 270.495
R435 VSS.n1936 VSS.n176 270.495
R436 VSS.n1937 VSS.n1936 270.495
R437 VSS.n1938 VSS.n1937 270.495
R438 VSS.n1938 VSS.n172 270.495
R439 VSS.n1945 VSS.n172 270.495
R440 VSS.n1946 VSS.n1945 270.495
R441 VSS.n1947 VSS.n1946 270.495
R442 VSS.n2185 VSS.n2184 263.776
R443 VSS.n1791 VSS.n1790 261.077
R444 VSS.n2372 VSS.n10 260.783
R445 VSS.n654 VSS.n650 253.755
R446 VSS.n2094 VSS.n2093 253.214
R447 VSS.n2093 VSS.n2092 253.214
R448 VSS.n2092 VSS.n2059 253.214
R449 VSS.n2086 VSS.n2059 253.214
R450 VSS.n2086 VSS.n2085 253.214
R451 VSS.n2085 VSS.n2084 253.214
R452 VSS.n2084 VSS.n2064 253.214
R453 VSS.n2078 VSS.n2064 253.214
R454 VSS.n2078 VSS.n2077 253.214
R455 VSS.n2077 VSS.n2076 253.214
R456 VSS.n2076 VSS.n2068 253.214
R457 VSS.n2070 VSS.n2068 253.214
R458 VSS.n10 VSS.n2 250.683
R459 VSS.n745 VSS.n744 250.536
R460 VSS.n358 VSS.n354 246.151
R461 VSS.n1378 VSS.n1256 246.151
R462 VSS.n447 VSS.n446 246.151
R463 VSS.n1201 VSS.n458 246.151
R464 VSS.n1947 VSS.n156 246.151
R465 VSS.n571 VSS.n542 242.81
R466 VSS.n572 VSS.n571 242.81
R467 VSS.n573 VSS.n572 242.81
R468 VSS.n573 VSS.n538 242.81
R469 VSS.n579 VSS.n538 242.81
R470 VSS.n580 VSS.n579 242.81
R471 VSS.n581 VSS.n580 242.81
R472 VSS.n587 VSS.n534 242.81
R473 VSS.n588 VSS.n587 242.81
R474 VSS.n589 VSS.n588 242.81
R475 VSS.n589 VSS.n530 242.81
R476 VSS.n595 VSS.n530 242.81
R477 VSS.n596 VSS.n595 242.81
R478 VSS.n598 VSS.n596 242.81
R479 VSS.n598 VSS.n597 242.81
R480 VSS.n632 VSS.n520 242.81
R481 VSS.n632 VSS.n523 242.81
R482 VSS.n739 VSS.n523 242.81
R483 VSS.n740 VSS.n739 239.167
R484 VSS.n2109 VSS.n2108 228.954
R485 VSS.n2110 VSS.n2109 228.954
R486 VSS.n2110 VSS.n103 228.954
R487 VSS.n2116 VSS.n103 228.954
R488 VSS.n2117 VSS.n2116 228.954
R489 VSS.n2118 VSS.n2117 228.954
R490 VSS.n2057 VSS.n118 213.608
R491 VSS.n886 VSS.n885 210.766
R492 VSS.n885 VSS.n884 210.766
R493 VSS.n884 VSS.n841 210.766
R494 VSS.n878 VSS.n841 210.766
R495 VSS.n878 VSS.n877 210.766
R496 VSS.n877 VSS.n876 210.766
R497 VSS.n876 VSS.n845 210.766
R498 VSS.n870 VSS.n869 210.766
R499 VSS.n869 VSS.n868 210.766
R500 VSS.n868 VSS.n850 210.766
R501 VSS.n862 VSS.n850 210.766
R502 VSS.n862 VSS.n861 210.766
R503 VSS.n861 VSS.n860 210.766
R504 VSS.n860 VSS.n854 210.766
R505 VSS.n854 VSS.n307 210.766
R506 VSS.n407 VSS.n405 210.766
R507 VSS.n407 VSS.n406 210.766
R508 VSS.n406 VSS.n327 210.766
R509 VSS.n953 VSS.n952 210.766
R510 VSS.n952 VSS.n951 210.766
R511 VSS.n951 VSS.n909 210.766
R512 VSS.n945 VSS.n909 210.766
R513 VSS.n945 VSS.n944 210.766
R514 VSS.n944 VSS.n943 210.766
R515 VSS.n943 VSS.n913 210.766
R516 VSS.n937 VSS.n936 210.766
R517 VSS.n936 VSS.n935 210.766
R518 VSS.n935 VSS.n917 210.766
R519 VSS.n929 VSS.n917 210.766
R520 VSS.n929 VSS.n928 210.766
R521 VSS.n928 VSS.n927 210.766
R522 VSS.n927 VSS.n921 210.766
R523 VSS.n921 VSS.n291 210.766
R524 VSS.n1337 VSS.n1336 210.766
R525 VSS.n1338 VSS.n1337 210.766
R526 VSS.n1338 VSS.n329 210.766
R527 VSS.n992 VSS.n991 210.766
R528 VSS.n991 VSS.n990 210.766
R529 VSS.n990 VSS.n976 210.766
R530 VSS.n984 VSS.n976 210.766
R531 VSS.n984 VSS.n983 210.766
R532 VSS.n983 VSS.n982 210.766
R533 VSS.n982 VSS.n268 210.766
R534 VSS.n1654 VSS.n269 210.766
R535 VSS.n1648 VSS.n269 210.766
R536 VSS.n1648 VSS.n1647 210.766
R537 VSS.n1647 VSS.n1646 210.766
R538 VSS.n1646 VSS.n275 210.766
R539 VSS.n1640 VSS.n275 210.766
R540 VSS.n1640 VSS.n1639 210.766
R541 VSS.n1639 VSS.n1638 210.766
R542 VSS.n336 VSS.n335 210.766
R543 VSS.n336 VSS.n331 210.766
R544 VSS.n1478 VSS.n331 210.766
R545 VSS.n1698 VSS.n255 210.766
R546 VSS.n1692 VSS.n255 210.766
R547 VSS.n1692 VSS.n1691 210.766
R548 VSS.n1691 VSS.n1690 210.766
R549 VSS.n1690 VSS.n263 210.766
R550 VSS.n1684 VSS.n263 210.766
R551 VSS.n1684 VSS.n1683 210.766
R552 VSS.n1681 VSS.n1656 210.766
R553 VSS.n1675 VSS.n1656 210.766
R554 VSS.n1675 VSS.n1674 210.766
R555 VSS.n1674 VSS.n1673 210.766
R556 VSS.n1673 VSS.n1660 210.766
R557 VSS.n1667 VSS.n1660 210.766
R558 VSS.n1667 VSS.n1666 210.766
R559 VSS.n1666 VSS.n1665 210.766
R560 VSS.n1905 VSS.n189 210.766
R561 VSS.n1911 VSS.n189 210.766
R562 VSS.n1912 VSS.n1911 210.766
R563 VSS.n2302 VSS.n2301 207.837
R564 VSS.n2054 VSS.n123 207.668
R565 VSS.n2048 VSS.n123 207.668
R566 VSS.n2048 VSS.n2047 207.668
R567 VSS.n2047 VSS.n2046 207.668
R568 VSS.n2046 VSS.n2035 207.668
R569 VSS.n2040 VSS.n2035 207.668
R570 VSS.n2040 VSS.n2039 207.668
R571 VSS.n2039 VSS.n92 207.668
R572 VSS.n2186 VSS.n92 207.668
R573 VSS.n2193 VSS.n85 207.668
R574 VSS.n2194 VSS.n2193 207.668
R575 VSS.n2195 VSS.n2194 207.668
R576 VSS.n2195 VSS.n79 207.668
R577 VSS.n1483 VSS.n327 207.605
R578 VSS.n1481 VSS.n329 207.605
R579 VSS.n1479 VSS.n1478 207.605
R580 VSS.n1913 VSS.n1912 207.605
R581 VSS.n2344 VSS.n27 200.476
R582 VSS.n2010 VSS.n145 196.203
R583 VSS.n1853 VSS.n207 194.62
R584 VSS.n26 VSS.n20 193.958
R585 VSS.n2002 VSS.n130 192.245
R586 VSS.n2231 VSS.n79 191.054
R587 VSS.n701 VSS.n700 172.887
R588 VSS.n2294 VSS.n60 172.149
R589 VSS.n1775 VSS.n118 170.887
R590 VSS.n1440 VSS.n1439 167.708
R591 VSS.n1377 VSS.n1257 167.708
R592 VSS.n1396 VSS.n1395 167.708
R593 VSS.n1211 VSS.n462 167.708
R594 VSS.n1957 VSS.n160 167.708
R595 VSS.n116 VSS.n107 163.702
R596 VSS.n2281 VSS.n71 162.431
R597 VSS.n2027 VSS.n131 158.228
R598 VSS.n2027 VSS.n2026 158.228
R599 VSS.n2058 VSS.n116 154.267
R600 VSS.n534 VSS.n518 150.542
R601 VSS.n2271 VSS.n78 138.831
R602 VSS.n2272 VSS.n2271 138.831
R603 VSS.n2353 VSS.n20 132.022
R604 VSS.n128 VSS.n122 131.869
R605 VSS.n2282 VSS.n2281 131.696
R606 VSS.n2384 VSS.n2383 131.672
R607 VSS.n545 VSS.n542 131.118
R608 VSS.n870 VSS.n849 130.674
R609 VSS.n937 VSS.n267 130.674
R610 VSS.n1655 VSS.n1654 130.674
R611 VSS.n1682 VSS.n1681 130.674
R612 VSS.n2055 VSS.n122 129.792
R613 VSS.n27 VSS.n26 125.502
R614 VSS.n2138 VSS.n2137 124.343
R615 VSS.n2108 VSS.n107 123.635
R616 VSS.n2281 VSS.n2280 115.23
R617 VSS.n886 VSS.n833 113.814
R618 VSS.n953 VSS.n901 113.814
R619 VSS.n992 VSS.n968 113.814
R620 VSS.n1699 VSS.n1698 113.814
R621 VSS.n753 VSS.n752 103.141
R622 VSS.n760 VSS.n508 103.141
R623 VSS.n759 VSS.n509 103.141
R624 VSS.n766 VSS.n504 103.141
R625 VSS.n768 VSS.n767 103.141
R626 VSS.n1161 VSS.n499 103.141
R627 VSS.n823 VSS.n492 103.141
R628 VSS.n1153 VSS.n1152 103.141
R629 VSS.n1136 VSS.n824 103.141
R630 VSS.n1146 VSS.n1137 103.141
R631 VSS.n1145 VSS.n1139 103.141
R632 VSS.n1138 VSS.n323 103.141
R633 VSS.n744 VSS.n519 101.981
R634 VSS.n2028 VSS.n128 99.9337
R635 VSS.t30 VSS.n117 95.2243
R636 VSS.n597 VSS.n519 93.482
R637 VSS.n581 VSS.n518 92.268
R638 VSS.n1523 VSS.n117 88.5219
R639 VSS.n1561 VSS.n117 88.5219
R640 VSS.n279 VSS.n117 88.5219
R641 VSS.n195 VSS.n117 88.5219
R642 VSS.n1808 VSS.n128 85.4435
R643 VSS.n1523 VSS.n307 81.1451
R644 VSS.n1561 VSS.n291 81.1451
R645 VSS.n1638 VSS.n279 81.1451
R646 VSS.n1665 VSS.n195 81.1451
R647 VSS.n849 VSS.n845 80.0913
R648 VSS.n913 VSS.n267 80.0913
R649 VSS.n1655 VSS.n268 80.0913
R650 VSS.n1683 VSS.n1682 80.0913
R651 VSS.n751 VSS.n513 77.9039
R652 VSS.n2055 VSS.n2054 77.8759
R653 VSS.n2139 VSS.n2138 77.8759
R654 VSS.n2303 VSS.n2302 75.3694
R655 VSS.n1486 VSS.n1485 75.1609
R656 VSS.n2138 VSS.n85 63.3392
R657 VSS.n1790 VSS.n1789 55.3802
R658 VSS.n1166 VSS.n1165 54.3135
R659 VSS.n2094 VSS.n2058 54.1874
R660 VSS.n1160 VSS.n490 52.6676
R661 VSS.n2185 VSS.n2139 51.9174
R662 VSS.n2186 VSS.n2185 47.7641
R663 VSS.n744 VSS.n520 47.3483
R664 VSS.n405 VSS.n117 41.0997
R665 VSS.n1336 VSS.n117 41.0997
R666 VSS.n335 VSS.n117 41.0997
R667 VSS.n1905 VSS.n117 41.0997
R668 VSS.n207 VSS.n128 36.3929
R669 VSS.n145 VSS.n138 28.4815
R670 VSS.n1485 VSS.n325 27.9799
R671 VSS.n742 VSS.n513 25.2368
R672 VSS.n701 VSS.n654 25.097
R673 VSS.n1440 VSS.n358 24.3451
R674 VSS.n1378 VSS.n1377 24.3451
R675 VSS.n1396 VSS.n447 24.3451
R676 VSS.n462 VSS.n458 24.3451
R677 VSS.n160 VSS.n156 24.3451
R678 VSS.n2057 VSS.n116 20.7673
R679 VSS.n702 VSS.n653 19.3426
R680 VSS.n2382 VSS.n6 18.4216
R681 VSS.n2378 VSS.n2377 18.4216
R682 VSS.n2374 VSS.n2373 18.4216
R683 VSS.n2373 VSS.n9 18.4216
R684 VSS.n2369 VSS.n9 18.4216
R685 VSS.n2369 VSS.n12 18.4216
R686 VSS.n2364 VSS.n12 18.4216
R687 VSS.n2364 VSS.n15 18.4216
R688 VSS.n2360 VSS.n15 18.4216
R689 VSS.n2360 VSS.n17 18.4216
R690 VSS.n2356 VSS.n17 18.4216
R691 VSS.n2356 VSS.n19 18.4216
R692 VSS.n2352 VSS.n19 18.4216
R693 VSS.n2352 VSS.n21 18.4216
R694 VSS.n2107 VSS.n106 18.4216
R695 VSS.n2111 VSS.n106 18.4216
R696 VSS.n2111 VSS.n104 18.4216
R697 VSS.n2115 VSS.n104 18.4216
R698 VSS.n2115 VSS.n102 18.4216
R699 VSS.n2119 VSS.n102 18.4216
R700 VSS.n2119 VSS.n99 18.4216
R701 VSS.n2136 VSS.n99 18.4216
R702 VSS.n2136 VSS.n100 18.4216
R703 VSS.n2132 VSS.n2131 18.4216
R704 VSS.n2128 VSS.n2127 18.4216
R705 VSS.n2124 VSS.n2123 18.4216
R706 VSS.n1906 VSS.n190 18.4216
R707 VSS.n1910 VSS.n190 18.4216
R708 VSS.n1910 VSS.n187 18.4216
R709 VSS.n1915 VSS.n187 18.4216
R710 VSS.n1915 VSS.n185 18.4216
R711 VSS.n1919 VSS.n185 18.4216
R712 VSS.n1919 VSS.n183 18.4216
R713 VSS.n1923 VSS.n183 18.4216
R714 VSS.n1923 VSS.n181 18.4216
R715 VSS.n1927 VSS.n181 18.4216
R716 VSS.n1927 VSS.n179 18.4216
R717 VSS.n1931 VSS.n179 18.4216
R718 VSS.n1931 VSS.n177 18.4216
R719 VSS.n1935 VSS.n177 18.4216
R720 VSS.n1935 VSS.n175 18.4216
R721 VSS.n1939 VSS.n175 18.4216
R722 VSS.n1939 VSS.n173 18.4216
R723 VSS.n1944 VSS.n173 18.4216
R724 VSS.n1944 VSS.n170 18.4216
R725 VSS.n1948 VSS.n170 18.4216
R726 VSS.n1949 VSS.n1948 18.4216
R727 VSS.n1697 VSS.n257 18.4216
R728 VSS.n1693 VSS.n257 18.4216
R729 VSS.n1693 VSS.n262 18.4216
R730 VSS.n1689 VSS.n262 18.4216
R731 VSS.n1689 VSS.n264 18.4216
R732 VSS.n1685 VSS.n264 18.4216
R733 VSS.n1685 VSS.n266 18.4216
R734 VSS.n1680 VSS.n266 18.4216
R735 VSS.n1680 VSS.n1657 18.4216
R736 VSS.n1676 VSS.n1657 18.4216
R737 VSS.n1676 VSS.n1659 18.4216
R738 VSS.n1672 VSS.n1659 18.4216
R739 VSS.n1672 VSS.n1661 18.4216
R740 VSS.n1668 VSS.n1661 18.4216
R741 VSS.n1668 VSS.n1664 18.4216
R742 VSS.n1664 VSS.n192 18.4216
R743 VSS.n993 VSS.n975 18.4216
R744 VSS.n989 VSS.n975 18.4216
R745 VSS.n989 VSS.n977 18.4216
R746 VSS.n985 VSS.n977 18.4216
R747 VSS.n985 VSS.n979 18.4216
R748 VSS.n981 VSS.n979 18.4216
R749 VSS.n981 VSS.n270 18.4216
R750 VSS.n1653 VSS.n270 18.4216
R751 VSS.n1653 VSS.n271 18.4216
R752 VSS.n1649 VSS.n271 18.4216
R753 VSS.n1649 VSS.n274 18.4216
R754 VSS.n1645 VSS.n274 18.4216
R755 VSS.n1645 VSS.n276 18.4216
R756 VSS.n1641 VSS.n276 18.4216
R757 VSS.n1641 VSS.n278 18.4216
R758 VSS.n1637 VSS.n278 18.4216
R759 VSS.n954 VSS.n908 18.4216
R760 VSS.n950 VSS.n908 18.4216
R761 VSS.n950 VSS.n910 18.4216
R762 VSS.n946 VSS.n910 18.4216
R763 VSS.n946 VSS.n912 18.4216
R764 VSS.n942 VSS.n912 18.4216
R765 VSS.n942 VSS.n914 18.4216
R766 VSS.n938 VSS.n914 18.4216
R767 VSS.n938 VSS.n916 18.4216
R768 VSS.n934 VSS.n916 18.4216
R769 VSS.n934 VSS.n918 18.4216
R770 VSS.n930 VSS.n918 18.4216
R771 VSS.n930 VSS.n920 18.4216
R772 VSS.n926 VSS.n920 18.4216
R773 VSS.n926 VSS.n922 18.4216
R774 VSS.n922 VSS.n300 18.4216
R775 VSS.n887 VSS.n840 18.4216
R776 VSS.n883 VSS.n840 18.4216
R777 VSS.n883 VSS.n842 18.4216
R778 VSS.n879 VSS.n842 18.4216
R779 VSS.n879 VSS.n844 18.4216
R780 VSS.n875 VSS.n844 18.4216
R781 VSS.n875 VSS.n846 18.4216
R782 VSS.n871 VSS.n846 18.4216
R783 VSS.n871 VSS.n848 18.4216
R784 VSS.n867 VSS.n848 18.4216
R785 VSS.n867 VSS.n851 18.4216
R786 VSS.n863 VSS.n851 18.4216
R787 VSS.n863 VSS.n853 18.4216
R788 VSS.n859 VSS.n853 18.4216
R789 VSS.n859 VSS.n855 18.4216
R790 VSS.n855 VSS.n316 18.4216
R791 VSS.n782 VSS.n780 18.4216
R792 VSS.n786 VSS.n779 18.4216
R793 VSS.n790 VSS.n788 18.4216
R794 VSS.n794 VSS.n777 18.4216
R795 VSS.n798 VSS.n796 18.4216
R796 VSS.n802 VSS.n775 18.4216
R797 VSS.n805 VSS.n804 18.4216
R798 VSS.n809 VSS.n808 18.4216
R799 VSS.n633 VSS.n631 18.4216
R800 VSS.n633 VSS.n524 18.4216
R801 VSS.n738 VSS.n524 18.4216
R802 VSS.n738 VSS.n525 18.4216
R803 VSS.n734 VSS.n525 18.4216
R804 VSS.n734 VSS.n637 18.4216
R805 VSS.n730 VSS.n637 18.4216
R806 VSS.n730 VSS.n639 18.4216
R807 VSS.n726 VSS.n639 18.4216
R808 VSS.n726 VSS.n641 18.4216
R809 VSS.n722 VSS.n641 18.4216
R810 VSS.n722 VSS.n643 18.4216
R811 VSS.n718 VSS.n643 18.4216
R812 VSS.n718 VSS.n645 18.4216
R813 VSS.n714 VSS.n645 18.4216
R814 VSS.n714 VSS.n647 18.4216
R815 VSS.n710 VSS.n647 18.4216
R816 VSS.n710 VSS.n649 18.4216
R817 VSS.n706 VSS.n649 18.4216
R818 VSS.n706 VSS.n651 18.4216
R819 VSS.n702 VSS.n651 18.4216
R820 VSS.n408 VSS.n317 18.4216
R821 VSS.n408 VSS.n403 18.4216
R822 VSS.n412 VSS.n403 18.4216
R823 VSS.n413 VSS.n412 18.4216
R824 VSS.n415 VSS.n413 18.4216
R825 VSS.n415 VSS.n401 18.4216
R826 VSS.n419 VSS.n401 18.4216
R827 VSS.n419 VSS.n399 18.4216
R828 VSS.n423 VSS.n399 18.4216
R829 VSS.n423 VSS.n397 18.4216
R830 VSS.n427 VSS.n397 18.4216
R831 VSS.n427 VSS.n395 18.4216
R832 VSS.n431 VSS.n395 18.4216
R833 VSS.n431 VSS.n393 18.4216
R834 VSS.n435 VSS.n393 18.4216
R835 VSS.n435 VSS.n391 18.4216
R836 VSS.n439 VSS.n391 18.4216
R837 VSS.n439 VSS.n389 18.4216
R838 VSS.n444 VSS.n389 18.4216
R839 VSS.n444 VSS.n387 18.4216
R840 VSS.n1397 VSS.n387 18.4216
R841 VSS.n337 VSS.n334 18.4216
R842 VSS.n337 VSS.n332 18.4216
R843 VSS.n1477 VSS.n332 18.4216
R844 VSS.n1477 VSS.n333 18.4216
R845 VSS.n1473 VSS.n333 18.4216
R846 VSS.n1473 VSS.n341 18.4216
R847 VSS.n1469 VSS.n341 18.4216
R848 VSS.n1469 VSS.n343 18.4216
R849 VSS.n1465 VSS.n343 18.4216
R850 VSS.n1465 VSS.n345 18.4216
R851 VSS.n1461 VSS.n345 18.4216
R852 VSS.n1461 VSS.n347 18.4216
R853 VSS.n1457 VSS.n347 18.4216
R854 VSS.n1457 VSS.n349 18.4216
R855 VSS.n1453 VSS.n349 18.4216
R856 VSS.n1453 VSS.n351 18.4216
R857 VSS.n1449 VSS.n351 18.4216
R858 VSS.n1449 VSS.n353 18.4216
R859 VSS.n1445 VSS.n353 18.4216
R860 VSS.n1445 VSS.n355 18.4216
R861 VSS.n1441 VSS.n355 18.4216
R862 VSS.n1335 VSS.n301 18.4216
R863 VSS.n1339 VSS.n1335 18.4216
R864 VSS.n1340 VSS.n1339 18.4216
R865 VSS.n1340 VSS.n1331 18.4216
R866 VSS.n1344 VSS.n1331 18.4216
R867 VSS.n1344 VSS.n1330 18.4216
R868 VSS.n1348 VSS.n1330 18.4216
R869 VSS.n1348 VSS.n1328 18.4216
R870 VSS.n1352 VSS.n1328 18.4216
R871 VSS.n1352 VSS.n1326 18.4216
R872 VSS.n1356 VSS.n1326 18.4216
R873 VSS.n1356 VSS.n1324 18.4216
R874 VSS.n1360 VSS.n1324 18.4216
R875 VSS.n1360 VSS.n1322 18.4216
R876 VSS.n1364 VSS.n1322 18.4216
R877 VSS.n1364 VSS.n1320 18.4216
R878 VSS.n1368 VSS.n1320 18.4216
R879 VSS.n1368 VSS.n1318 18.4216
R880 VSS.n1372 VSS.n1318 18.4216
R881 VSS.n1372 VSS.n1258 18.4216
R882 VSS.n1376 VSS.n1258 18.4216
R883 VSS.n817 VSS.n816 18.4216
R884 VSS.n1169 VSS.n489 18.4216
R885 VSS.n1169 VSS.n487 18.4216
R886 VSS.n1173 VSS.n487 18.4216
R887 VSS.n1173 VSS.n485 18.4216
R888 VSS.n1177 VSS.n485 18.4216
R889 VSS.n1177 VSS.n483 18.4216
R890 VSS.n1181 VSS.n483 18.4216
R891 VSS.n1181 VSS.n481 18.4216
R892 VSS.n1185 VSS.n481 18.4216
R893 VSS.n1185 VSS.n479 18.4216
R894 VSS.n1189 VSS.n479 18.4216
R895 VSS.n1189 VSS.n477 18.4216
R896 VSS.n1193 VSS.n477 18.4216
R897 VSS.n1193 VSS.n475 18.4216
R898 VSS.n1198 VSS.n475 18.4216
R899 VSS.n1198 VSS.n472 18.4216
R900 VSS.n1202 VSS.n472 18.4216
R901 VSS.n1203 VSS.n1202 18.4216
R902 VSS.n570 VSS.n543 18.4216
R903 VSS.n570 VSS.n541 18.4216
R904 VSS.n574 VSS.n541 18.4216
R905 VSS.n574 VSS.n539 18.4216
R906 VSS.n578 VSS.n539 18.4216
R907 VSS.n578 VSS.n537 18.4216
R908 VSS.n582 VSS.n537 18.4216
R909 VSS.n582 VSS.n535 18.4216
R910 VSS.n586 VSS.n535 18.4216
R911 VSS.n586 VSS.n533 18.4216
R912 VSS.n590 VSS.n533 18.4216
R913 VSS.n590 VSS.n531 18.4216
R914 VSS.n594 VSS.n531 18.4216
R915 VSS.n594 VSS.n529 18.4216
R916 VSS.n599 VSS.n529 18.4216
R917 VSS.n599 VSS.n527 18.4216
R918 VSS.n564 VSS.n563 18.4216
R919 VSS.n561 VSS.n547 18.4216
R920 VSS.n557 VSS.n556 18.4216
R921 VSS.n554 VSS.n551 18.4216
R922 VSS.n551 VSS.n516 18.4216
R923 VSS.n746 VSS.n516 18.4216
R924 VSS.n746 VSS.n514 18.4216
R925 VSS.n750 VSS.n514 18.4216
R926 VSS.n750 VSS.n507 18.4216
R927 VSS.n761 VSS.n507 18.4216
R928 VSS.n761 VSS.n505 18.4216
R929 VSS.n765 VSS.n505 18.4216
R930 VSS.n765 VSS.n498 18.4216
R931 VSS.n1162 VSS.n498 18.4216
R932 VSS.n1164 VSS.n494 18.4216
R933 VSS.n1151 VSS.n494 18.4216
R934 VSS.n1151 VSS.n825 18.4216
R935 VSS.n1147 VSS.n825 18.4216
R936 VSS.n1147 VSS.n1135 18.4216
R937 VSS.n1135 VSS.n1134 18.4216
R938 VSS.n1134 VSS.n827 18.4216
R939 VSS.n1130 VSS.n827 18.4216
R940 VSS.n1130 VSS.n829 18.4216
R941 VSS.n1127 VSS.n830 18.4216
R942 VSS.n1123 VSS.n1122 18.4216
R943 VSS.n1120 VSS.n834 18.4216
R944 VSS.n1116 VSS.n1115 18.4216
R945 VSS.n1107 VSS.n890 18.4216
R946 VSS.n1103 VSS.n1102 18.4216
R947 VSS.n1100 VSS.n893 18.4216
R948 VSS.n1096 VSS.n1095 18.4216
R949 VSS.n1095 VSS.n896 18.4216
R950 VSS.n1092 VSS.n897 18.4216
R951 VSS.n1088 VSS.n1087 18.4216
R952 VSS.n1085 VSS.n902 18.4216
R953 VSS.n1081 VSS.n1080 18.4216
R954 VSS.n1072 VSS.n957 18.4216
R955 VSS.n1068 VSS.n1067 18.4216
R956 VSS.n1065 VSS.n960 18.4216
R957 VSS.n1061 VSS.n1060 18.4216
R958 VSS.n1060 VSS.n963 18.4216
R959 VSS.n1057 VSS.n964 18.4216
R960 VSS.n1053 VSS.n1052 18.4216
R961 VSS.n1050 VSS.n969 18.4216
R962 VSS.n1046 VSS.n1045 18.4216
R963 VSS.n1037 VSS.n996 18.4216
R964 VSS.n1033 VSS.n1032 18.4216
R965 VSS.n1030 VSS.n999 18.4216
R966 VSS.n1026 VSS.n1025 18.4216
R967 VSS.n1025 VSS.n1002 18.4216
R968 VSS.n1022 VSS.n1003 18.4216
R969 VSS.n1018 VSS.n1017 18.4216
R970 VSS.n1014 VSS.n1013 18.4216
R971 VSS.n1010 VSS.n1009 18.4216
R972 VSS.n248 VSS.n247 18.4216
R973 VSS.n253 VSS.n241 18.4216
R974 VSS.n1702 VSS.n1701 18.4216
R975 VSS.n1706 VSS.n1705 18.4216
R976 VSS.n1709 VSS.n1706 18.4216
R977 VSS.n1713 VSS.n237 18.4216
R978 VSS.n1717 VSS.n1715 18.4216
R979 VSS.n1721 VSS.n235 18.4216
R980 VSS.n1724 VSS.n1723 18.4216
R981 VSS.n1771 VSS.n1730 18.4216
R982 VSS.n1767 VSS.n1766 18.4216
R983 VSS.n1762 VSS.n1761 18.4216
R984 VSS.n1758 VSS.n1757 18.4216
R985 VSS.n1754 VSS.n1753 18.4216
R986 VSS.n1753 VSS.n1752 18.4216
R987 VSS.n1750 VSS.n1734 18.4216
R988 VSS.n1746 VSS.n1745 18.4216
R989 VSS.n1743 VSS.n1739 18.4216
R990 VSS.n2103 VSS.n2102 18.4216
R991 VSS.n2100 VSS.n112 18.4216
R992 VSS.n2096 VSS.n2095 18.4216
R993 VSS.n2095 VSS.n115 18.4216
R994 VSS.n2091 VSS.n115 18.4216
R995 VSS.n2091 VSS.n2060 18.4216
R996 VSS.n2087 VSS.n2060 18.4216
R997 VSS.n2087 VSS.n2063 18.4216
R998 VSS.n2083 VSS.n2063 18.4216
R999 VSS.n2083 VSS.n2065 18.4216
R1000 VSS.n2079 VSS.n2065 18.4216
R1001 VSS.n2079 VSS.n2067 18.4216
R1002 VSS.n2075 VSS.n2067 18.4216
R1003 VSS.n2075 VSS.n2069 18.4216
R1004 VSS.n2071 VSS.n2069 18.4216
R1005 VSS.n2071 VSS.n5 18.4216
R1006 VSS.n1776 VSS.n230 18.4216
R1007 VSS.n1780 VSS.n230 18.4216
R1008 VSS.n1780 VSS.n228 18.4216
R1009 VSS.n1784 VSS.n228 18.4216
R1010 VSS.n1784 VSS.n226 18.4216
R1011 VSS.n1788 VSS.n226 18.4216
R1012 VSS.n1788 VSS.n221 18.4216
R1013 VSS.n1793 VSS.n221 18.4216
R1014 VSS.n1793 VSS.n219 18.4216
R1015 VSS.n1797 VSS.n219 18.4216
R1016 VSS.n1797 VSS.n217 18.4216
R1017 VSS.n1801 VSS.n217 18.4216
R1018 VSS.n1801 VSS.n215 18.4216
R1019 VSS.n1805 VSS.n215 18.4216
R1020 VSS.n1805 VSS.n213 18.4216
R1021 VSS.n1809 VSS.n213 18.4216
R1022 VSS.n1854 VSS.n1812 18.4216
R1023 VSS.n1850 VSS.n1812 18.4216
R1024 VSS.n1850 VSS.n1814 18.4216
R1025 VSS.n1846 VSS.n1814 18.4216
R1026 VSS.n1846 VSS.n1816 18.4216
R1027 VSS.n1842 VSS.n1816 18.4216
R1028 VSS.n1842 VSS.n1818 18.4216
R1029 VSS.n1838 VSS.n1818 18.4216
R1030 VSS.n1838 VSS.n1820 18.4216
R1031 VSS.n1834 VSS.n1820 18.4216
R1032 VSS.n1834 VSS.n1822 18.4216
R1033 VSS.n1830 VSS.n1822 18.4216
R1034 VSS.n1830 VSS.n1824 18.4216
R1035 VSS.n1826 VSS.n1824 18.4216
R1036 VSS.n1826 VSS.n133 18.4216
R1037 VSS.n2025 VSS.n133 18.4216
R1038 VSS.n2025 VSS.n134 18.4216
R1039 VSS.n2021 VSS.n134 18.4216
R1040 VSS.n2021 VSS.n137 18.4216
R1041 VSS.n2017 VSS.n137 18.4216
R1042 VSS.n2017 VSS.n139 18.4216
R1043 VSS.n627 VSS.n604 18.4216
R1044 VSS.n623 VSS.n622 18.4216
R1045 VSS.n620 VSS.n607 18.4216
R1046 VSS.n616 VSS.n615 18.4216
R1047 VSS.n615 VSS.n614 18.4216
R1048 VSS.n612 VSS.n512 18.4216
R1049 VSS.n754 VSS.n512 18.4216
R1050 VSS.n754 VSS.n510 18.4216
R1051 VSS.n758 VSS.n510 18.4216
R1052 VSS.n758 VSS.n503 18.4216
R1053 VSS.n769 VSS.n503 18.4216
R1054 VSS.n769 VSS.n500 18.4216
R1055 VSS.n1159 VSS.n500 18.4216
R1056 VSS.n1155 VSS.n1154 18.4216
R1057 VSS.n1154 VSS.n822 18.4216
R1058 VSS.n1140 VSS.n822 18.4216
R1059 VSS.n1144 VSS.n1140 18.4216
R1060 VSS.n1144 VSS.n322 18.4216
R1061 VSS.n1487 VSS.n322 18.4216
R1062 VSS.n1487 VSS.n320 18.4216
R1063 VSS.n1492 VSS.n320 18.4216
R1064 VSS.n1492 VSS.n319 18.4216
R1065 VSS.n1496 VSS.n1495 18.4216
R1066 VSS.n1500 VSS.n1499 18.4216
R1067 VSS.n1504 VSS.n1503 18.4216
R1068 VSS.n1508 VSS.n1507 18.4216
R1069 VSS.n1517 VSS.n1516 18.4216
R1070 VSS.n1521 VSS.n314 18.4216
R1071 VSS.n1525 VSS.n306 18.4216
R1072 VSS.n1530 VSS.n304 18.4216
R1073 VSS.n1530 VSS.n303 18.4216
R1074 VSS.n1534 VSS.n1533 18.4216
R1075 VSS.n1538 VSS.n1537 18.4216
R1076 VSS.n1542 VSS.n1541 18.4216
R1077 VSS.n1546 VSS.n1545 18.4216
R1078 VSS.n1555 VSS.n1554 18.4216
R1079 VSS.n1559 VSS.n298 18.4216
R1080 VSS.n1563 VSS.n290 18.4216
R1081 VSS.n1568 VSS.n288 18.4216
R1082 VSS.n1568 VSS.n287 18.4216
R1083 VSS.n1573 VSS.n1571 18.4216
R1084 VSS.n1577 VSS.n285 18.4216
R1085 VSS.n1580 VSS.n1579 18.4216
R1086 VSS.n1584 VSS.n1583 18.4216
R1087 VSS.n1631 VSS.n1630 18.4216
R1088 VSS.n1628 VSS.n1590 18.4216
R1089 VSS.n1624 VSS.n1623 18.4216
R1090 VSS.n1621 VSS.n1593 18.4216
R1091 VSS.n1617 VSS.n1593 18.4216
R1092 VSS.n1615 VSS.n1614 18.4216
R1093 VSS.n1612 VSS.n1597 18.4216
R1094 VSS.n1608 VSS.n1607 18.4216
R1095 VSS.n1605 VSS.n1601 18.4216
R1096 VSS.n1901 VSS.n196 18.4216
R1097 VSS.n1897 VSS.n1896 18.4216
R1098 VSS.n1894 VSS.n199 18.4216
R1099 VSS.n1890 VSS.n1889 18.4216
R1100 VSS.n1889 VSS.n202 18.4216
R1101 VSS.n1886 VSS.n203 18.4216
R1102 VSS.n1882 VSS.n1881 18.4216
R1103 VSS.n1879 VSS.n208 18.4216
R1104 VSS.n1875 VSS.n1874 18.4216
R1105 VSS.n1866 VSS.n1865 18.4216
R1106 VSS.n1863 VSS.n1858 18.4216
R1107 VSS.n1859 VSS.n127 18.4216
R1108 VSS.n2030 VSS.n124 18.4216
R1109 VSS.n2053 VSS.n124 18.4216
R1110 VSS.n2053 VSS.n125 18.4216
R1111 VSS.n2049 VSS.n125 18.4216
R1112 VSS.n2049 VSS.n2034 18.4216
R1113 VSS.n2045 VSS.n2034 18.4216
R1114 VSS.n2045 VSS.n2036 18.4216
R1115 VSS.n2041 VSS.n2036 18.4216
R1116 VSS.n2041 VSS.n2038 18.4216
R1117 VSS.n2038 VSS.n90 18.4216
R1118 VSS.n2187 VSS.n90 18.4216
R1119 VSS.n2192 VSS.n86 18.4216
R1120 VSS.n2192 VSS.n84 18.4216
R1121 VSS.n2196 VSS.n84 18.4216
R1122 VSS.n2196 VSS.n81 18.4216
R1123 VSS.n2229 VSS.n81 18.4216
R1124 VSS.n2229 VSS.n82 18.4216
R1125 VSS.n2225 VSS.n82 18.4216
R1126 VSS.n2225 VSS.n2200 18.4216
R1127 VSS.n2221 VSS.n2200 18.4216
R1128 VSS.n2221 VSS.n2202 18.4216
R1129 VSS.n2217 VSS.n2202 18.4216
R1130 VSS.n2217 VSS.n2215 18.4216
R1131 VSS.n2215 VSS.n2214 18.4216
R1132 VSS.n2212 VSS.n2205 18.4216
R1133 VSS.n2208 VSS.n2207 18.4216
R1134 VSS.n2345 VSS.n25 18.4216
R1135 VSS.n2341 VSS.n25 18.4216
R1136 VSS.n2341 VSS.n29 18.4216
R1137 VSS.n2337 VSS.n29 18.4216
R1138 VSS.n2337 VSS.n32 18.4216
R1139 VSS.n2333 VSS.n32 18.4216
R1140 VSS.n2333 VSS.n34 18.4216
R1141 VSS.n2329 VSS.n34 18.4216
R1142 VSS.n2329 VSS.n36 18.4216
R1143 VSS.n2325 VSS.n36 18.4216
R1144 VSS.n2325 VSS.n38 18.4216
R1145 VSS.n2321 VSS.n38 18.4216
R1146 VSS.n2321 VSS.n40 18.4216
R1147 VSS.n2317 VSS.n40 18.4216
R1148 VSS.n2317 VSS.n42 18.4216
R1149 VSS.n2313 VSS.n42 18.4216
R1150 VSS.n2313 VSS.n44 18.4216
R1151 VSS.n2309 VSS.n44 18.4216
R1152 VSS.n2309 VSS.n46 18.4216
R1153 VSS.n2305 VSS.n46 18.4216
R1154 VSS.n2305 VSS.n48 18.4216
R1155 VSS.n661 VSS.n660 18.4216
R1156 VSS.n663 VSS.n657 18.4216
R1157 VSS.n698 VSS.n658 18.4216
R1158 VSS.n694 VSS.n658 18.4216
R1159 VSS.n694 VSS.n669 18.4216
R1160 VSS.n690 VSS.n669 18.4216
R1161 VSS.n690 VSS.n672 18.4216
R1162 VSS.n686 VSS.n672 18.4216
R1163 VSS.n686 VSS.n683 18.4216
R1164 VSS.n683 VSS.n682 18.4216
R1165 VSS.n679 VSS.n678 18.4216
R1166 VSS.n675 VSS.n674 18.4216
R1167 VSS.n1209 VSS.n467 18.4216
R1168 VSS.n1213 VSS.n461 18.4216
R1169 VSS.n1217 VSS.n459 18.4216
R1170 VSS.n1217 VSS.n457 18.4216
R1171 VSS.n1221 VSS.n457 18.4216
R1172 VSS.n1221 VSS.n454 18.4216
R1173 VSS.n1226 VSS.n454 18.4216
R1174 VSS.n1226 VSS.n452 18.4216
R1175 VSS.n1230 VSS.n452 18.4216
R1176 VSS.n1231 VSS.n1230 18.4216
R1177 VSS.n1233 VSS.n449 18.4216
R1178 VSS.n1237 VSS.n450 18.4216
R1179 VSS.n1244 VSS.n1243 18.4216
R1180 VSS.n1246 VSS.n1241 18.4216
R1181 VSS.n1393 VSS.n1242 18.4216
R1182 VSS.n1389 VSS.n1242 18.4216
R1183 VSS.n1389 VSS.n1249 18.4216
R1184 VSS.n1385 VSS.n1249 18.4216
R1185 VSS.n1385 VSS.n1252 18.4216
R1186 VSS.n1381 VSS.n1252 18.4216
R1187 VSS.n1381 VSS.n1254 18.4216
R1188 VSS.n1262 VSS.n1254 18.4216
R1189 VSS.n1266 VSS.n1264 18.4216
R1190 VSS.n1270 VSS.n1259 18.4216
R1191 VSS.n1313 VSS.n1273 18.4216
R1192 VSS.n1309 VSS.n1308 18.4216
R1193 VSS.n1306 VSS.n1276 18.4216
R1194 VSS.n1302 VSS.n1276 18.4216
R1195 VSS.n1302 VSS.n1277 18.4216
R1196 VSS.n1298 VSS.n1277 18.4216
R1197 VSS.n1298 VSS.n1279 18.4216
R1198 VSS.n1294 VSS.n1279 18.4216
R1199 VSS.n1294 VSS.n1291 18.4216
R1200 VSS.n1291 VSS.n1290 18.4216
R1201 VSS.n1287 VSS.n1286 18.4216
R1202 VSS.n1283 VSS.n1282 18.4216
R1203 VSS.n370 VSS.n369 18.4216
R1204 VSS.n372 VSS.n366 18.4216
R1205 VSS.n1437 VSS.n367 18.4216
R1206 VSS.n1433 VSS.n367 18.4216
R1207 VSS.n1433 VSS.n1408 18.4216
R1208 VSS.n1429 VSS.n1408 18.4216
R1209 VSS.n1429 VSS.n1411 18.4216
R1210 VSS.n1425 VSS.n1411 18.4216
R1211 VSS.n1425 VSS.n1422 18.4216
R1212 VSS.n1422 VSS.n1421 18.4216
R1213 VSS.n1418 VSS.n1417 18.4216
R1214 VSS.n1414 VSS.n1413 18.4216
R1215 VSS.n1955 VSS.n165 18.4216
R1216 VSS.n1959 VSS.n159 18.4216
R1217 VSS.n1963 VSS.n157 18.4216
R1218 VSS.n1963 VSS.n155 18.4216
R1219 VSS.n1967 VSS.n155 18.4216
R1220 VSS.n1967 VSS.n151 18.4216
R1221 VSS.n1972 VSS.n151 18.4216
R1222 VSS.n1972 VSS.n149 18.4216
R1223 VSS.n1976 VSS.n149 18.4216
R1224 VSS.n1977 VSS.n1976 18.4216
R1225 VSS.n1979 VSS.n147 18.4216
R1226 VSS.n1983 VSS.n144 18.4216
R1227 VSS.n1987 VSS.n1986 18.4216
R1228 VSS.n2008 VSS.n1988 18.4216
R1229 VSS.n2004 VSS.n2003 18.4216
R1230 VSS.n2003 VSS.n1992 18.4216
R1231 VSS.n1999 VSS.n1992 18.4216
R1232 VSS.n1999 VSS.n1994 18.4216
R1233 VSS.n1994 VSS.n69 18.4216
R1234 VSS.n2284 VSS.n69 18.4216
R1235 VSS.n2284 VSS.n66 18.4216
R1236 VSS.n2293 VSS.n66 18.4216
R1237 VSS.n2293 VSS.n67 18.4216
R1238 VSS.n2289 VSS.n2288 18.4216
R1239 VSS.n2295 VSS.n58 18.4216
R1240 VSS.n62 VSS.n57 18.4216
R1241 VSS.n2237 VSS.n2236 18.4216
R1242 VSS.n2239 VSS.n2232 18.4216
R1243 VSS.n2268 VSS.n2232 18.4216
R1244 VSS.n2268 VSS.n2234 18.4216
R1245 VSS.n2264 VSS.n2234 18.4216
R1246 VSS.n2264 VSS.n2243 18.4216
R1247 VSS.n2260 VSS.n2243 18.4216
R1248 VSS.n2260 VSS.n2245 18.4216
R1249 VSS.n2256 VSS.n2245 18.4216
R1250 VSS.n2256 VSS.n2253 18.4216
R1251 VSS.n2253 VSS.n2252 18.4216
R1252 VSS.n2252 VSS.n2247 18.4216
R1253 VSS.n2248 VSS.n51 18.4216
R1254 VSS.n2150 VSS.n2148 18.4216
R1255 VSS.n2154 VSS.n2144 18.4216
R1256 VSS.n2158 VSS.n2156 18.4216
R1257 VSS.n2183 VSS.n2141 18.4216
R1258 VSS.n2183 VSS.n2142 18.4216
R1259 VSS.n2179 VSS.n2142 18.4216
R1260 VSS.n2179 VSS.n2162 18.4216
R1261 VSS.n2175 VSS.n2162 18.4216
R1262 VSS.n2175 VSS.n2164 18.4216
R1263 VSS.n2166 VSS.n2164 18.4216
R1264 VSS.n2170 VSS.n2166 18.4216
R1265 VSS.n2170 VSS.n77 18.4216
R1266 VSS.n2274 VSS.n77 18.4216
R1267 VSS.n2274 VSS.n73 18.4216
R1268 VSS.n2279 VSS.n73 18.4216
R1269 VSS.n2279 VSS.n75 18.4216
R1270 VSS.n75 VSS.n74 18.4216
R1271 VSS.n566 VSS.n543 17.8689
R1272 VSS.n2299 VSS.n48 17.8689
R1273 VSS.n2382 VSS.n5 16.3952
R1274 VSS.n630 VSS.n629 12.5268
R1275 VSS.n1155 VSS.n501 12.5268
R1276 VSS.n1513 VSS.n1512 12.5268
R1277 VSS.n1551 VSS.n1550 12.5268
R1278 VSS.n1633 VSS.n280 12.5268
R1279 VSS.n1904 VSS.n1903 12.5268
R1280 VSS.n1868 VSS.n211 12.5268
R1281 VSS.n91 VSS.n86 12.5268
R1282 VSS.n456 VSS.t25 12.3005
R1283 VSS.n376 VSS.t19 12.3005
R1284 VSS.n1996 VSS.t21 12.3005
R1285 VSS.n153 VSS.t29 12.3005
R1286 VSS.n375 VSS.t23 12.3005
R1287 VSS.n379 VSS.t17 12.3005
R1288 VSS.n666 VSS.t27 12.3005
R1289 VSS.n1164 VSS.n493 11.4216
R1290 VSS.n1109 VSS.n837 11.4216
R1291 VSS.n1074 VSS.n905 11.4216
R1292 VSS.n1039 VSS.n972 11.4216
R1293 VSS.n258 VSS.n256 11.4216
R1294 VSS.n1774 VSS.n1773 11.4216
R1295 VSS.n2103 VSS.n108 11.4216
R1296 VSS.n1204 VSS.n470 11.4216
R1297 VSS.n1398 VSS.n385 11.4216
R1298 VSS.n1316 VSS.n1315 11.4216
R1299 VSS.n363 VSS.n357 11.4216
R1300 VSS.n1950 VSS.n168 11.4216
R1301 VSS.n2012 VSS.n142 11.4216
R1302 VSS.n59 VSS.n57 11.4216
R1303 VSS.n0 VSS.t34 11.2214
R1304 VSS.n744 VSS.n743 10.9728
R1305 VSS.n324 VSS.n117 10.9728
R1306 VSS.n2385 VSS.n2384 10.4005
R1307 VSS.n2384 VSS.n0 10.4005
R1308 VSS.n1162 VSS.n493 9.94787
R1309 VSS.n1113 VSS.n837 9.94787
R1310 VSS.n1078 VSS.n905 9.94787
R1311 VSS.n1043 VSS.n972 9.94787
R1312 VSS.n1005 VSS.n256 9.94787
R1313 VSS.n1774 VSS.n1728 9.94787
R1314 VSS.n1737 VSS.n108 9.94787
R1315 VSS.n1205 VSS.n1204 9.94787
R1316 VSS.n1399 VSS.n1398 9.94787
R1317 VSS.n1316 VSS.n1272 9.94787
R1318 VSS.n361 VSS.n357 9.94787
R1319 VSS.n1951 VSS.n1950 9.94787
R1320 VSS.n2013 VSS.n2012 9.94787
R1321 VSS.n2295 VSS.n59 9.94787
R1322 VSS.n1159 VSS.n501 8.84261
R1323 VSS.n1512 VSS.n1511 8.84261
R1324 VSS.n1550 VSS.n1549 8.84261
R1325 VSS.n1586 VSS.n280 8.84261
R1326 VSS.n1904 VSS.n193 8.84261
R1327 VSS.n1872 VSS.n211 8.84261
R1328 VSS.n2187 VSS.n91 8.84261
R1329 VSS.n2347 VSS.n2346 8.84261
R1330 VSS.n1167 VSS.n1166 8.77835
R1331 VSS.n1950 VSS.n1949 7.92155
R1332 VSS.n1398 VSS.n1397 7.92155
R1333 VSS.n1441 VSS.n357 7.92155
R1334 VSS.n1376 VSS.n1316 7.92155
R1335 VSS.n1204 VSS.n1203 7.92155
R1336 VSS.n2012 VSS.n139 7.92155
R1337 VSS.n74 VSS.n59 7.92155
R1338 VSS.n1906 VSS.n1904 7.82945
R1339 VSS.n631 VSS.n630 7.82945
R1340 VSS.n1512 VSS.n317 7.82945
R1341 VSS.n334 VSS.n280 7.82945
R1342 VSS.n1550 VSS.n301 7.82945
R1343 VSS.n819 VSS.n501 7.82945
R1344 VSS.n1854 VSS.n211 7.82945
R1345 VSS.n2346 VSS.n2345 7.82945
R1346 VSS.n2146 VSS.n91 7.82945
R1347 VSS.n743 VSS.n742 6.58389
R1348 VSS.n753 VSS.n751 6.58389
R1349 VSS.n752 VSS.n508 6.58389
R1350 VSS.n760 VSS.n759 6.58389
R1351 VSS.n509 VSS.n504 6.58389
R1352 VSS.n768 VSS.n766 6.58389
R1353 VSS.n767 VSS.n499 6.58389
R1354 VSS.n1161 VSS.n1160 6.58389
R1355 VSS.n1165 VSS.n492 6.58389
R1356 VSS.n1153 VSS.n823 6.58389
R1357 VSS.n1152 VSS.n824 6.58389
R1358 VSS.n1137 VSS.n1136 6.58389
R1359 VSS.n1146 VSS.n1145 6.58389
R1360 VSS.n1139 VSS.n1138 6.58389
R1361 VSS.n1486 VSS.n323 6.58389
R1362 VSS.n325 VSS.n324 6.58389
R1363 VSS.n2107 VSS.n108 6.44787
R1364 VSS.n1697 VSS.n256 6.44787
R1365 VSS.n993 VSS.n972 6.44787
R1366 VSS.n954 VSS.n905 6.44787
R1367 VSS.n887 VSS.n837 6.44787
R1368 VSS.n780 VSS.n493 6.44787
R1369 VSS.n1776 VSS.n1774 6.44787
R1370 VSS.n1166 VSS.n491 6.05199
R1371 VSS.n1442 VSS.n1441 5.2005
R1372 VSS.n1441 VSS.n1440 5.2005
R1373 VSS.n1443 VSS.n355 5.2005
R1374 VSS.n355 VSS.n354 5.2005
R1375 VSS.n1445 VSS.n1444 5.2005
R1376 VSS.n1446 VSS.n1445 5.2005
R1377 VSS.n353 VSS.n352 5.2005
R1378 VSS.n1447 VSS.n353 5.2005
R1379 VSS.n1450 VSS.n1449 5.2005
R1380 VSS.n1449 VSS.n1448 5.2005
R1381 VSS.n1451 VSS.n351 5.2005
R1382 VSS.n351 VSS.n350 5.2005
R1383 VSS.n1453 VSS.n1452 5.2005
R1384 VSS.n1454 VSS.n1453 5.2005
R1385 VSS.n349 VSS.n348 5.2005
R1386 VSS.n1455 VSS.n349 5.2005
R1387 VSS.n1458 VSS.n1457 5.2005
R1388 VSS.n1457 VSS.n1456 5.2005
R1389 VSS.n1459 VSS.n347 5.2005
R1390 VSS.n347 VSS.n346 5.2005
R1391 VSS.n1461 VSS.n1460 5.2005
R1392 VSS.n1462 VSS.n1461 5.2005
R1393 VSS.n345 VSS.n344 5.2005
R1394 VSS.n1463 VSS.n345 5.2005
R1395 VSS.n1466 VSS.n1465 5.2005
R1396 VSS.n1465 VSS.n1464 5.2005
R1397 VSS.n1467 VSS.n343 5.2005
R1398 VSS.n343 VSS.n342 5.2005
R1399 VSS.n1469 VSS.n1468 5.2005
R1400 VSS.n1470 VSS.n1469 5.2005
R1401 VSS.n341 VSS.n340 5.2005
R1402 VSS.n1471 VSS.n341 5.2005
R1403 VSS.n1474 VSS.n1473 5.2005
R1404 VSS.n1473 VSS.n1472 5.2005
R1405 VSS.n1475 VSS.n333 5.2005
R1406 VSS.n333 VSS.n330 5.2005
R1407 VSS.n1376 VSS.n1375 5.2005
R1408 VSS.n1377 VSS.n1376 5.2005
R1409 VSS.n1374 VSS.n1258 5.2005
R1410 VSS.n1258 VSS.n1256 5.2005
R1411 VSS.n1373 VSS.n1372 5.2005
R1412 VSS.n1372 VSS.n1371 5.2005
R1413 VSS.n1318 VSS.n1317 5.2005
R1414 VSS.n1370 VSS.n1318 5.2005
R1415 VSS.n1368 VSS.n1367 5.2005
R1416 VSS.n1369 VSS.n1368 5.2005
R1417 VSS.n1366 VSS.n1320 5.2005
R1418 VSS.n1320 VSS.n1319 5.2005
R1419 VSS.n1365 VSS.n1364 5.2005
R1420 VSS.n1364 VSS.n1363 5.2005
R1421 VSS.n1322 VSS.n1321 5.2005
R1422 VSS.n1362 VSS.n1322 5.2005
R1423 VSS.n1360 VSS.n1359 5.2005
R1424 VSS.n1361 VSS.n1360 5.2005
R1425 VSS.n1358 VSS.n1324 5.2005
R1426 VSS.n1324 VSS.n1323 5.2005
R1427 VSS.n1357 VSS.n1356 5.2005
R1428 VSS.n1356 VSS.n1355 5.2005
R1429 VSS.n1326 VSS.n1325 5.2005
R1430 VSS.n1354 VSS.n1326 5.2005
R1431 VSS.n1352 VSS.n1351 5.2005
R1432 VSS.n1353 VSS.n1352 5.2005
R1433 VSS.n1350 VSS.n1328 5.2005
R1434 VSS.n1328 VSS.n1327 5.2005
R1435 VSS.n1349 VSS.n1348 5.2005
R1436 VSS.n1348 VSS.n1347 5.2005
R1437 VSS.n1330 VSS.n1329 5.2005
R1438 VSS.n1346 VSS.n1330 5.2005
R1439 VSS.n1344 VSS.n1343 5.2005
R1440 VSS.n1345 VSS.n1344 5.2005
R1441 VSS.n1342 VSS.n1331 5.2005
R1442 VSS.n1331 VSS.n328 5.2005
R1443 VSS.n1397 VSS.n384 5.2005
R1444 VSS.n1397 VSS.n1396 5.2005
R1445 VSS.n442 VSS.n387 5.2005
R1446 VSS.n446 VSS.n387 5.2005
R1447 VSS.n444 VSS.n443 5.2005
R1448 VSS.n445 VSS.n444 5.2005
R1449 VSS.n441 VSS.n389 5.2005
R1450 VSS.n389 VSS.n388 5.2005
R1451 VSS.n440 VSS.n439 5.2005
R1452 VSS.n439 VSS.n438 5.2005
R1453 VSS.n391 VSS.n390 5.2005
R1454 VSS.n437 VSS.n391 5.2005
R1455 VSS.n435 VSS.n434 5.2005
R1456 VSS.n436 VSS.n435 5.2005
R1457 VSS.n433 VSS.n393 5.2005
R1458 VSS.n393 VSS.n392 5.2005
R1459 VSS.n432 VSS.n431 5.2005
R1460 VSS.n431 VSS.n430 5.2005
R1461 VSS.n395 VSS.n394 5.2005
R1462 VSS.n429 VSS.n395 5.2005
R1463 VSS.n427 VSS.n426 5.2005
R1464 VSS.n428 VSS.n427 5.2005
R1465 VSS.n425 VSS.n397 5.2005
R1466 VSS.n397 VSS.n396 5.2005
R1467 VSS.n424 VSS.n423 5.2005
R1468 VSS.n423 VSS.n422 5.2005
R1469 VSS.n399 VSS.n398 5.2005
R1470 VSS.n421 VSS.n399 5.2005
R1471 VSS.n419 VSS.n418 5.2005
R1472 VSS.n420 VSS.n419 5.2005
R1473 VSS.n417 VSS.n401 5.2005
R1474 VSS.n401 VSS.n400 5.2005
R1475 VSS.n416 VSS.n415 5.2005
R1476 VSS.n415 VSS.n414 5.2005
R1477 VSS.n413 VSS.n402 5.2005
R1478 VSS.n413 VSS.n326 5.2005
R1479 VSS.n1203 VSS.n469 5.2005
R1480 VSS.n1203 VSS.n462 5.2005
R1481 VSS.n1202 VSS.n473 5.2005
R1482 VSS.n1202 VSS.n1201 5.2005
R1483 VSS.n1196 VSS.n472 5.2005
R1484 VSS.n1200 VSS.n472 5.2005
R1485 VSS.n1198 VSS.n1197 5.2005
R1486 VSS.n1199 VSS.n1198 5.2005
R1487 VSS.n1195 VSS.n475 5.2005
R1488 VSS.n475 VSS.n474 5.2005
R1489 VSS.n1194 VSS.n1193 5.2005
R1490 VSS.n1193 VSS.n1192 5.2005
R1491 VSS.n477 VSS.n476 5.2005
R1492 VSS.n1191 VSS.n477 5.2005
R1493 VSS.n1189 VSS.n1188 5.2005
R1494 VSS.n1190 VSS.n1189 5.2005
R1495 VSS.n1187 VSS.n479 5.2005
R1496 VSS.n479 VSS.n478 5.2005
R1497 VSS.n1186 VSS.n1185 5.2005
R1498 VSS.n1185 VSS.n1184 5.2005
R1499 VSS.n481 VSS.n480 5.2005
R1500 VSS.n1183 VSS.n481 5.2005
R1501 VSS.n1181 VSS.n1180 5.2005
R1502 VSS.n1182 VSS.n1181 5.2005
R1503 VSS.n1179 VSS.n483 5.2005
R1504 VSS.n483 VSS.n482 5.2005
R1505 VSS.n1178 VSS.n1177 5.2005
R1506 VSS.n1177 VSS.n1176 5.2005
R1507 VSS.n485 VSS.n484 5.2005
R1508 VSS.n1175 VSS.n485 5.2005
R1509 VSS.n1173 VSS.n1172 5.2005
R1510 VSS.n1174 VSS.n1173 5.2005
R1511 VSS.n1171 VSS.n487 5.2005
R1512 VSS.n487 VSS.n486 5.2005
R1513 VSS.n1170 VSS.n1169 5.2005
R1514 VSS.n1169 VSS.n1168 5.2005
R1515 VSS.n736 VSS.n525 5.2005
R1516 VSS.n525 VSS.n522 5.2005
R1517 VSS.n735 VSS.n734 5.2005
R1518 VSS.n734 VSS.n733 5.2005
R1519 VSS.n637 VSS.n636 5.2005
R1520 VSS.n732 VSS.n637 5.2005
R1521 VSS.n730 VSS.n729 5.2005
R1522 VSS.n731 VSS.n730 5.2005
R1523 VSS.n728 VSS.n639 5.2005
R1524 VSS.n639 VSS.n638 5.2005
R1525 VSS.n727 VSS.n726 5.2005
R1526 VSS.n726 VSS.n725 5.2005
R1527 VSS.n641 VSS.n640 5.2005
R1528 VSS.n724 VSS.n641 5.2005
R1529 VSS.n722 VSS.n721 5.2005
R1530 VSS.n723 VSS.n722 5.2005
R1531 VSS.n720 VSS.n643 5.2005
R1532 VSS.n643 VSS.n642 5.2005
R1533 VSS.n719 VSS.n718 5.2005
R1534 VSS.n718 VSS.n717 5.2005
R1535 VSS.n645 VSS.n644 5.2005
R1536 VSS.n716 VSS.n645 5.2005
R1537 VSS.n714 VSS.n713 5.2005
R1538 VSS.n715 VSS.n714 5.2005
R1539 VSS.n712 VSS.n647 5.2005
R1540 VSS.n647 VSS.n646 5.2005
R1541 VSS.n711 VSS.n710 5.2005
R1542 VSS.n710 VSS.n709 5.2005
R1543 VSS.n649 VSS.n648 5.2005
R1544 VSS.n708 VSS.n649 5.2005
R1545 VSS.n706 VSS.n705 5.2005
R1546 VSS.n707 VSS.n706 5.2005
R1547 VSS.n704 VSS.n651 5.2005
R1548 VSS.n651 VSS.n650 5.2005
R1549 VSS.n703 VSS.n702 5.2005
R1550 VSS.n702 VSS.n701 5.2005
R1551 VSS.n631 VSS.n526 5.2005
R1552 VSS.n631 VSS.n520 5.2005
R1553 VSS.n634 VSS.n633 5.2005
R1554 VSS.n633 VSS.n632 5.2005
R1555 VSS.n635 VSS.n524 5.2005
R1556 VSS.n524 VSS.n523 5.2005
R1557 VSS.n738 VSS.n737 5.2005
R1558 VSS.n739 VSS.n738 5.2005
R1559 VSS.n812 VSS.n811 5.2005
R1560 VSS.n809 VSS.n772 5.2005
R1561 VSS.n808 VSS.n807 5.2005
R1562 VSS.n806 VSS.n805 5.2005
R1563 VSS.n804 VSS.n774 5.2005
R1564 VSS.n802 VSS.n801 5.2005
R1565 VSS.n800 VSS.n775 5.2005
R1566 VSS.n799 VSS.n798 5.2005
R1567 VSS.n796 VSS.n776 5.2005
R1568 VSS.n794 VSS.n793 5.2005
R1569 VSS.n792 VSS.n777 5.2005
R1570 VSS.n791 VSS.n790 5.2005
R1571 VSS.n788 VSS.n778 5.2005
R1572 VSS.n786 VSS.n785 5.2005
R1573 VSS.n784 VSS.n779 5.2005
R1574 VSS.n783 VSS.n782 5.2005
R1575 VSS.n780 VSS.n497 5.2005
R1576 VSS.n780 VSS.n490 5.2005
R1577 VSS.n489 VSS.n488 5.2005
R1578 VSS.n816 VSS.n815 5.2005
R1579 VSS.n817 VSS.n813 5.2005
R1580 VSS.n820 VSS.n819 5.2005
R1581 VSS.n856 VSS.n316 5.2005
R1582 VSS.n316 VSS.n307 5.2005
R1583 VSS.n857 VSS.n855 5.2005
R1584 VSS.n855 VSS.n854 5.2005
R1585 VSS.n859 VSS.n858 5.2005
R1586 VSS.n860 VSS.n859 5.2005
R1587 VSS.n853 VSS.n852 5.2005
R1588 VSS.n861 VSS.n853 5.2005
R1589 VSS.n864 VSS.n863 5.2005
R1590 VSS.n863 VSS.n862 5.2005
R1591 VSS.n865 VSS.n851 5.2005
R1592 VSS.n851 VSS.n850 5.2005
R1593 VSS.n867 VSS.n866 5.2005
R1594 VSS.n868 VSS.n867 5.2005
R1595 VSS.n848 VSS.n847 5.2005
R1596 VSS.n869 VSS.n848 5.2005
R1597 VSS.n872 VSS.n871 5.2005
R1598 VSS.n871 VSS.n870 5.2005
R1599 VSS.n873 VSS.n846 5.2005
R1600 VSS.n846 VSS.n845 5.2005
R1601 VSS.n875 VSS.n874 5.2005
R1602 VSS.n876 VSS.n875 5.2005
R1603 VSS.n844 VSS.n843 5.2005
R1604 VSS.n877 VSS.n844 5.2005
R1605 VSS.n880 VSS.n879 5.2005
R1606 VSS.n879 VSS.n878 5.2005
R1607 VSS.n881 VSS.n842 5.2005
R1608 VSS.n842 VSS.n841 5.2005
R1609 VSS.n883 VSS.n882 5.2005
R1610 VSS.n884 VSS.n883 5.2005
R1611 VSS.n840 VSS.n839 5.2005
R1612 VSS.n885 VSS.n840 5.2005
R1613 VSS.n888 VSS.n887 5.2005
R1614 VSS.n887 VSS.n886 5.2005
R1615 VSS.n412 VSS.n411 5.2005
R1616 VSS.n412 VSS.n327 5.2005
R1617 VSS.n410 VSS.n403 5.2005
R1618 VSS.n406 VSS.n403 5.2005
R1619 VSS.n409 VSS.n408 5.2005
R1620 VSS.n408 VSS.n407 5.2005
R1621 VSS.n404 VSS.n317 5.2005
R1622 VSS.n405 VSS.n317 5.2005
R1623 VSS.n923 VSS.n300 5.2005
R1624 VSS.n300 VSS.n291 5.2005
R1625 VSS.n924 VSS.n922 5.2005
R1626 VSS.n922 VSS.n921 5.2005
R1627 VSS.n926 VSS.n925 5.2005
R1628 VSS.n927 VSS.n926 5.2005
R1629 VSS.n920 VSS.n919 5.2005
R1630 VSS.n928 VSS.n920 5.2005
R1631 VSS.n931 VSS.n930 5.2005
R1632 VSS.n930 VSS.n929 5.2005
R1633 VSS.n932 VSS.n918 5.2005
R1634 VSS.n918 VSS.n917 5.2005
R1635 VSS.n934 VSS.n933 5.2005
R1636 VSS.n935 VSS.n934 5.2005
R1637 VSS.n916 VSS.n915 5.2005
R1638 VSS.n936 VSS.n916 5.2005
R1639 VSS.n939 VSS.n938 5.2005
R1640 VSS.n938 VSS.n937 5.2005
R1641 VSS.n940 VSS.n914 5.2005
R1642 VSS.n914 VSS.n913 5.2005
R1643 VSS.n942 VSS.n941 5.2005
R1644 VSS.n943 VSS.n942 5.2005
R1645 VSS.n912 VSS.n911 5.2005
R1646 VSS.n944 VSS.n912 5.2005
R1647 VSS.n947 VSS.n946 5.2005
R1648 VSS.n946 VSS.n945 5.2005
R1649 VSS.n948 VSS.n910 5.2005
R1650 VSS.n910 VSS.n909 5.2005
R1651 VSS.n950 VSS.n949 5.2005
R1652 VSS.n951 VSS.n950 5.2005
R1653 VSS.n908 VSS.n907 5.2005
R1654 VSS.n952 VSS.n908 5.2005
R1655 VSS.n955 VSS.n954 5.2005
R1656 VSS.n954 VSS.n953 5.2005
R1657 VSS.n1341 VSS.n1340 5.2005
R1658 VSS.n1340 VSS.n329 5.2005
R1659 VSS.n1339 VSS.n1332 5.2005
R1660 VSS.n1339 VSS.n1338 5.2005
R1661 VSS.n1335 VSS.n1334 5.2005
R1662 VSS.n1337 VSS.n1335 5.2005
R1663 VSS.n1333 VSS.n301 5.2005
R1664 VSS.n1336 VSS.n301 5.2005
R1665 VSS.n1637 VSS.n1636 5.2005
R1666 VSS.n1638 VSS.n1637 5.2005
R1667 VSS.n278 VSS.n277 5.2005
R1668 VSS.n1639 VSS.n278 5.2005
R1669 VSS.n1642 VSS.n1641 5.2005
R1670 VSS.n1641 VSS.n1640 5.2005
R1671 VSS.n1643 VSS.n276 5.2005
R1672 VSS.n276 VSS.n275 5.2005
R1673 VSS.n1645 VSS.n1644 5.2005
R1674 VSS.n1646 VSS.n1645 5.2005
R1675 VSS.n274 VSS.n273 5.2005
R1676 VSS.n1647 VSS.n274 5.2005
R1677 VSS.n1650 VSS.n1649 5.2005
R1678 VSS.n1649 VSS.n1648 5.2005
R1679 VSS.n1651 VSS.n271 5.2005
R1680 VSS.n271 VSS.n269 5.2005
R1681 VSS.n1653 VSS.n1652 5.2005
R1682 VSS.n1654 VSS.n1653 5.2005
R1683 VSS.n272 VSS.n270 5.2005
R1684 VSS.n270 VSS.n268 5.2005
R1685 VSS.n981 VSS.n980 5.2005
R1686 VSS.n982 VSS.n981 5.2005
R1687 VSS.n979 VSS.n978 5.2005
R1688 VSS.n983 VSS.n979 5.2005
R1689 VSS.n986 VSS.n985 5.2005
R1690 VSS.n985 VSS.n984 5.2005
R1691 VSS.n987 VSS.n977 5.2005
R1692 VSS.n977 VSS.n976 5.2005
R1693 VSS.n989 VSS.n988 5.2005
R1694 VSS.n990 VSS.n989 5.2005
R1695 VSS.n975 VSS.n974 5.2005
R1696 VSS.n991 VSS.n975 5.2005
R1697 VSS.n994 VSS.n993 5.2005
R1698 VSS.n993 VSS.n992 5.2005
R1699 VSS.n1477 VSS.n1476 5.2005
R1700 VSS.n1478 VSS.n1477 5.2005
R1701 VSS.n339 VSS.n332 5.2005
R1702 VSS.n332 VSS.n331 5.2005
R1703 VSS.n338 VSS.n337 5.2005
R1704 VSS.n337 VSS.n336 5.2005
R1705 VSS.n334 VSS.n281 5.2005
R1706 VSS.n335 VSS.n334 5.2005
R1707 VSS.n1662 VSS.n192 5.2005
R1708 VSS.n1665 VSS.n192 5.2005
R1709 VSS.n1664 VSS.n1663 5.2005
R1710 VSS.n1666 VSS.n1664 5.2005
R1711 VSS.n1669 VSS.n1668 5.2005
R1712 VSS.n1668 VSS.n1667 5.2005
R1713 VSS.n1670 VSS.n1661 5.2005
R1714 VSS.n1661 VSS.n1660 5.2005
R1715 VSS.n1672 VSS.n1671 5.2005
R1716 VSS.n1673 VSS.n1672 5.2005
R1717 VSS.n1659 VSS.n1658 5.2005
R1718 VSS.n1674 VSS.n1659 5.2005
R1719 VSS.n1677 VSS.n1676 5.2005
R1720 VSS.n1676 VSS.n1675 5.2005
R1721 VSS.n1678 VSS.n1657 5.2005
R1722 VSS.n1657 VSS.n1656 5.2005
R1723 VSS.n1680 VSS.n1679 5.2005
R1724 VSS.n1681 VSS.n1680 5.2005
R1725 VSS.n266 VSS.n265 5.2005
R1726 VSS.n1683 VSS.n266 5.2005
R1727 VSS.n1686 VSS.n1685 5.2005
R1728 VSS.n1685 VSS.n1684 5.2005
R1729 VSS.n1687 VSS.n264 5.2005
R1730 VSS.n264 VSS.n263 5.2005
R1731 VSS.n1689 VSS.n1688 5.2005
R1732 VSS.n1690 VSS.n1689 5.2005
R1733 VSS.n262 VSS.n261 5.2005
R1734 VSS.n1691 VSS.n262 5.2005
R1735 VSS.n1694 VSS.n1693 5.2005
R1736 VSS.n1693 VSS.n1692 5.2005
R1737 VSS.n1695 VSS.n257 5.2005
R1738 VSS.n257 VSS.n255 5.2005
R1739 VSS.n1697 VSS.n1696 5.2005
R1740 VSS.n1698 VSS.n1697 5.2005
R1741 VSS.n187 VSS.n186 5.2005
R1742 VSS.n1912 VSS.n187 5.2005
R1743 VSS.n1910 VSS.n1909 5.2005
R1744 VSS.n1911 VSS.n1910 5.2005
R1745 VSS.n1908 VSS.n190 5.2005
R1746 VSS.n190 VSS.n189 5.2005
R1747 VSS.n1907 VSS.n1906 5.2005
R1748 VSS.n1906 VSS.n1905 5.2005
R1749 VSS.n1949 VSS.n167 5.2005
R1750 VSS.n1949 VSS.n160 5.2005
R1751 VSS.n1948 VSS.n171 5.2005
R1752 VSS.n1948 VSS.n1947 5.2005
R1753 VSS.n1942 VSS.n170 5.2005
R1754 VSS.n1946 VSS.n170 5.2005
R1755 VSS.n1944 VSS.n1943 5.2005
R1756 VSS.n1945 VSS.n1944 5.2005
R1757 VSS.n1941 VSS.n173 5.2005
R1758 VSS.n173 VSS.n172 5.2005
R1759 VSS.n1940 VSS.n1939 5.2005
R1760 VSS.n1939 VSS.n1938 5.2005
R1761 VSS.n175 VSS.n174 5.2005
R1762 VSS.n1937 VSS.n175 5.2005
R1763 VSS.n1935 VSS.n1934 5.2005
R1764 VSS.n1936 VSS.n1935 5.2005
R1765 VSS.n1933 VSS.n177 5.2005
R1766 VSS.n177 VSS.n176 5.2005
R1767 VSS.n1932 VSS.n1931 5.2005
R1768 VSS.n1931 VSS.n1930 5.2005
R1769 VSS.n179 VSS.n178 5.2005
R1770 VSS.n1929 VSS.n179 5.2005
R1771 VSS.n1927 VSS.n1926 5.2005
R1772 VSS.n1928 VSS.n1927 5.2005
R1773 VSS.n1925 VSS.n181 5.2005
R1774 VSS.n181 VSS.n180 5.2005
R1775 VSS.n1924 VSS.n1923 5.2005
R1776 VSS.n1923 VSS.n1922 5.2005
R1777 VSS.n183 VSS.n182 5.2005
R1778 VSS.n1921 VSS.n183 5.2005
R1779 VSS.n1919 VSS.n1918 5.2005
R1780 VSS.n1920 VSS.n1919 5.2005
R1781 VSS.n1917 VSS.n185 5.2005
R1782 VSS.n185 VSS.n184 5.2005
R1783 VSS.n1916 VSS.n1915 5.2005
R1784 VSS.n1915 VSS.n1914 5.2005
R1785 VSS.n2120 VSS.n2119 5.2005
R1786 VSS.n2119 VSS.n2118 5.2005
R1787 VSS.n102 VSS.n101 5.2005
R1788 VSS.n2117 VSS.n102 5.2005
R1789 VSS.n2115 VSS.n2114 5.2005
R1790 VSS.n2116 VSS.n2115 5.2005
R1791 VSS.n2113 VSS.n104 5.2005
R1792 VSS.n104 VSS.n103 5.2005
R1793 VSS.n2112 VSS.n2111 5.2005
R1794 VSS.n2111 VSS.n2110 5.2005
R1795 VSS.n106 VSS.n105 5.2005
R1796 VSS.n2109 VSS.n106 5.2005
R1797 VSS.n2107 VSS.n2106 5.2005
R1798 VSS.n2108 VSS.n2107 5.2005
R1799 VSS.n2136 VSS.n2135 5.2005
R1800 VSS.n2137 VSS.n2136 5.2005
R1801 VSS.n2121 VSS.n99 5.2005
R1802 VSS.n99 VSS.n98 5.2005
R1803 VSS.n96 VSS.n88 5.2005
R1804 VSS.n2123 VSS.n2122 5.2005
R1805 VSS.n2125 VSS.n2124 5.2005
R1806 VSS.n2127 VSS.n2126 5.2005
R1807 VSS.n2129 VSS.n2128 5.2005
R1808 VSS.n2131 VSS.n2130 5.2005
R1809 VSS.n2133 VSS.n2132 5.2005
R1810 VSS.n2134 VSS.n100 5.2005
R1811 VSS.n2369 VSS.n2368 5.2005
R1812 VSS.n2370 VSS.n2369 5.2005
R1813 VSS.n13 VSS.n9 5.2005
R1814 VSS.n2371 VSS.n9 5.2005
R1815 VSS.n2373 VSS.n8 5.2005
R1816 VSS.n2373 VSS.n2372 5.2005
R1817 VSS.n2375 VSS.n2374 5.2005
R1818 VSS.n2377 VSS.n2376 5.2005
R1819 VSS.n2379 VSS.n2378 5.2005
R1820 VSS.n2380 VSS.n6 5.2005
R1821 VSS.n2382 VSS.n2381 5.2005
R1822 VSS.n2383 VSS.n2382 5.2005
R1823 VSS.n2350 VSS.n21 5.2005
R1824 VSS.n26 VSS.n21 5.2005
R1825 VSS.n2352 VSS.n2351 5.2005
R1826 VSS.n2353 VSS.n2352 5.2005
R1827 VSS.n19 VSS.n18 5.2005
R1828 VSS.n2354 VSS.n19 5.2005
R1829 VSS.n2357 VSS.n2356 5.2005
R1830 VSS.n2356 VSS.n2355 5.2005
R1831 VSS.n2358 VSS.n17 5.2005
R1832 VSS.n17 VSS.n16 5.2005
R1833 VSS.n2360 VSS.n2359 5.2005
R1834 VSS.n2361 VSS.n2360 5.2005
R1835 VSS.n15 VSS.n14 5.2005
R1836 VSS.n2362 VSS.n15 5.2005
R1837 VSS.n2365 VSS.n2364 5.2005
R1838 VSS.n2364 VSS.n2363 5.2005
R1839 VSS.n2366 VSS.n12 5.2005
R1840 VSS.n12 VSS.n11 5.2005
R1841 VSS.n568 VSS.n543 5.2005
R1842 VSS.n543 VSS.n542 5.2005
R1843 VSS.n570 VSS.n569 5.2005
R1844 VSS.n571 VSS.n570 5.2005
R1845 VSS.n541 VSS.n540 5.2005
R1846 VSS.n572 VSS.n541 5.2005
R1847 VSS.n575 VSS.n574 5.2005
R1848 VSS.n574 VSS.n573 5.2005
R1849 VSS.n576 VSS.n539 5.2005
R1850 VSS.n539 VSS.n538 5.2005
R1851 VSS.n578 VSS.n577 5.2005
R1852 VSS.n579 VSS.n578 5.2005
R1853 VSS.n537 VSS.n536 5.2005
R1854 VSS.n580 VSS.n537 5.2005
R1855 VSS.n583 VSS.n582 5.2005
R1856 VSS.n582 VSS.n581 5.2005
R1857 VSS.n584 VSS.n535 5.2005
R1858 VSS.n535 VSS.n534 5.2005
R1859 VSS.n586 VSS.n585 5.2005
R1860 VSS.n587 VSS.n586 5.2005
R1861 VSS.n533 VSS.n532 5.2005
R1862 VSS.n588 VSS.n533 5.2005
R1863 VSS.n591 VSS.n590 5.2005
R1864 VSS.n590 VSS.n589 5.2005
R1865 VSS.n592 VSS.n531 5.2005
R1866 VSS.n531 VSS.n530 5.2005
R1867 VSS.n594 VSS.n593 5.2005
R1868 VSS.n595 VSS.n594 5.2005
R1869 VSS.n529 VSS.n528 5.2005
R1870 VSS.n596 VSS.n529 5.2005
R1871 VSS.n600 VSS.n599 5.2005
R1872 VSS.n599 VSS.n598 5.2005
R1873 VSS.n601 VSS.n527 5.2005
R1874 VSS.n597 VSS.n527 5.2005
R1875 VSS.n7 VSS.n5 5.2005
R1876 VSS.n5 VSS.n2 5.2005
R1877 VSS.n2072 VSS.n2071 5.2005
R1878 VSS.n2071 VSS.n2070 5.2005
R1879 VSS.n2073 VSS.n2069 5.2005
R1880 VSS.n2069 VSS.n2068 5.2005
R1881 VSS.n2075 VSS.n2074 5.2005
R1882 VSS.n2076 VSS.n2075 5.2005
R1883 VSS.n2067 VSS.n2066 5.2005
R1884 VSS.n2077 VSS.n2067 5.2005
R1885 VSS.n2080 VSS.n2079 5.2005
R1886 VSS.n2079 VSS.n2078 5.2005
R1887 VSS.n2081 VSS.n2065 5.2005
R1888 VSS.n2065 VSS.n2064 5.2005
R1889 VSS.n2083 VSS.n2082 5.2005
R1890 VSS.n2084 VSS.n2083 5.2005
R1891 VSS.n2063 VSS.n2062 5.2005
R1892 VSS.n2085 VSS.n2063 5.2005
R1893 VSS.n2088 VSS.n2087 5.2005
R1894 VSS.n2087 VSS.n2086 5.2005
R1895 VSS.n2089 VSS.n2060 5.2005
R1896 VSS.n2060 VSS.n2059 5.2005
R1897 VSS.n2091 VSS.n2090 5.2005
R1898 VSS.n2092 VSS.n2091 5.2005
R1899 VSS.n2061 VSS.n115 5.2005
R1900 VSS.n2093 VSS.n115 5.2005
R1901 VSS.n2095 VSS.n113 5.2005
R1902 VSS.n2095 VSS.n2094 5.2005
R1903 VSS.n2097 VSS.n2096 5.2005
R1904 VSS.n2098 VSS.n112 5.2005
R1905 VSS.n2100 VSS.n2099 5.2005
R1906 VSS.n2102 VSS.n111 5.2005
R1907 VSS.n2104 VSS.n2103 5.2005
R1908 VSS.n2103 VSS.n107 5.2005
R1909 VSS.n1737 VSS.n109 5.2005
R1910 VSS.n1741 VSS.n1739 5.2005
R1911 VSS.n1743 VSS.n1742 5.2005
R1912 VSS.n1745 VSS.n1735 5.2005
R1913 VSS.n1747 VSS.n1746 5.2005
R1914 VSS.n1748 VSS.n1734 5.2005
R1915 VSS.n1750 VSS.n1749 5.2005
R1916 VSS.n1752 VSS.n1733 5.2005
R1917 VSS.n1753 VSS.n1732 5.2005
R1918 VSS.n1753 VSS.n107 5.2005
R1919 VSS.n1755 VSS.n1754 5.2005
R1920 VSS.n1757 VSS.n1756 5.2005
R1921 VSS.n1759 VSS.n1758 5.2005
R1922 VSS.n1761 VSS.n1760 5.2005
R1923 VSS.n1763 VSS.n1762 5.2005
R1924 VSS.n1766 VSS.n1764 5.2005
R1925 VSS.n1768 VSS.n1767 5.2005
R1926 VSS.n1769 VSS.n1730 5.2005
R1927 VSS.n1771 VSS.n1770 5.2005
R1928 VSS.n1773 VSS.n1729 5.2005
R1929 VSS.n1728 VSS.n1727 5.2005
R1930 VSS.n1725 VSS.n1724 5.2005
R1931 VSS.n1723 VSS.n234 5.2005
R1932 VSS.n1721 VSS.n1720 5.2005
R1933 VSS.n1719 VSS.n235 5.2005
R1934 VSS.n1718 VSS.n1717 5.2005
R1935 VSS.n1715 VSS.n236 5.2005
R1936 VSS.n1713 VSS.n1712 5.2005
R1937 VSS.n1711 VSS.n237 5.2005
R1938 VSS.n1710 VSS.n1709 5.2005
R1939 VSS.n1706 VSS.n238 5.2005
R1940 VSS.n1707 VSS.n1706 5.2005
R1941 VSS.n1705 VSS.n1704 5.2005
R1942 VSS.n1703 VSS.n1702 5.2005
R1943 VSS.n1701 VSS.n240 5.2005
R1944 VSS.n251 VSS.n241 5.2005
R1945 VSS.n253 VSS.n252 5.2005
R1946 VSS.n250 VSS.n247 5.2005
R1947 VSS.n249 VSS.n248 5.2005
R1948 VSS.n259 VSS.n258 5.2005
R1949 VSS.n1006 VSS.n1005 5.2005
R1950 VSS.n1009 VSS.n1008 5.2005
R1951 VSS.n1011 VSS.n1010 5.2005
R1952 VSS.n1013 VSS.n1012 5.2005
R1953 VSS.n1015 VSS.n1014 5.2005
R1954 VSS.n1017 VSS.n1016 5.2005
R1955 VSS.n1019 VSS.n1018 5.2005
R1956 VSS.n1020 VSS.n1003 5.2005
R1957 VSS.n1022 VSS.n1021 5.2005
R1958 VSS.n1004 VSS.n1002 5.2005
R1959 VSS.n1025 VSS.n1000 5.2005
R1960 VSS.n1025 VSS.n1024 5.2005
R1961 VSS.n1027 VSS.n1026 5.2005
R1962 VSS.n1028 VSS.n999 5.2005
R1963 VSS.n1030 VSS.n1029 5.2005
R1964 VSS.n1032 VSS.n997 5.2005
R1965 VSS.n1034 VSS.n1033 5.2005
R1966 VSS.n1035 VSS.n996 5.2005
R1967 VSS.n1037 VSS.n1036 5.2005
R1968 VSS.n1040 VSS.n1039 5.2005
R1969 VSS.n1043 VSS.n1042 5.2005
R1970 VSS.n1045 VSS.n970 5.2005
R1971 VSS.n1047 VSS.n1046 5.2005
R1972 VSS.n1048 VSS.n969 5.2005
R1973 VSS.n1050 VSS.n1049 5.2005
R1974 VSS.n1052 VSS.n966 5.2005
R1975 VSS.n1054 VSS.n1053 5.2005
R1976 VSS.n1055 VSS.n964 5.2005
R1977 VSS.n1057 VSS.n1056 5.2005
R1978 VSS.n965 VSS.n963 5.2005
R1979 VSS.n1060 VSS.n961 5.2005
R1980 VSS.n1060 VSS.n1059 5.2005
R1981 VSS.n1062 VSS.n1061 5.2005
R1982 VSS.n1063 VSS.n960 5.2005
R1983 VSS.n1065 VSS.n1064 5.2005
R1984 VSS.n1067 VSS.n958 5.2005
R1985 VSS.n1069 VSS.n1068 5.2005
R1986 VSS.n1070 VSS.n957 5.2005
R1987 VSS.n1072 VSS.n1071 5.2005
R1988 VSS.n1075 VSS.n1074 5.2005
R1989 VSS.n1078 VSS.n1077 5.2005
R1990 VSS.n1080 VSS.n903 5.2005
R1991 VSS.n1082 VSS.n1081 5.2005
R1992 VSS.n1083 VSS.n902 5.2005
R1993 VSS.n1085 VSS.n1084 5.2005
R1994 VSS.n1087 VSS.n899 5.2005
R1995 VSS.n1089 VSS.n1088 5.2005
R1996 VSS.n1090 VSS.n897 5.2005
R1997 VSS.n1092 VSS.n1091 5.2005
R1998 VSS.n898 VSS.n896 5.2005
R1999 VSS.n1095 VSS.n894 5.2005
R2000 VSS.n1095 VSS.n1094 5.2005
R2001 VSS.n1097 VSS.n1096 5.2005
R2002 VSS.n1098 VSS.n893 5.2005
R2003 VSS.n1100 VSS.n1099 5.2005
R2004 VSS.n1102 VSS.n891 5.2005
R2005 VSS.n1104 VSS.n1103 5.2005
R2006 VSS.n1105 VSS.n890 5.2005
R2007 VSS.n1107 VSS.n1106 5.2005
R2008 VSS.n1110 VSS.n1109 5.2005
R2009 VSS.n1113 VSS.n1112 5.2005
R2010 VSS.n1115 VSS.n835 5.2005
R2011 VSS.n1117 VSS.n1116 5.2005
R2012 VSS.n1118 VSS.n834 5.2005
R2013 VSS.n1120 VSS.n1119 5.2005
R2014 VSS.n1122 VSS.n831 5.2005
R2015 VSS.n1124 VSS.n1123 5.2005
R2016 VSS.n1125 VSS.n830 5.2005
R2017 VSS.n1127 VSS.n1126 5.2005
R2018 VSS.n829 VSS.n828 5.2005
R2019 VSS.n1131 VSS.n1130 5.2005
R2020 VSS.n1130 VSS.n1129 5.2005
R2021 VSS.n1132 VSS.n827 5.2005
R2022 VSS.n827 VSS.n325 5.2005
R2023 VSS.n1134 VSS.n1133 5.2005
R2024 VSS.n1134 VSS.n323 5.2005
R2025 VSS.n1135 VSS.n826 5.2005
R2026 VSS.n1139 VSS.n1135 5.2005
R2027 VSS.n1148 VSS.n1147 5.2005
R2028 VSS.n1147 VSS.n1146 5.2005
R2029 VSS.n1149 VSS.n825 5.2005
R2030 VSS.n1136 VSS.n825 5.2005
R2031 VSS.n1151 VSS.n1150 5.2005
R2032 VSS.n1152 VSS.n1151 5.2005
R2033 VSS.n496 VSS.n494 5.2005
R2034 VSS.n823 VSS.n494 5.2005
R2035 VSS.n1164 VSS.n1163 5.2005
R2036 VSS.n1165 VSS.n1164 5.2005
R2037 VSS.n1163 VSS.n1162 5.2005
R2038 VSS.n1162 VSS.n1161 5.2005
R2039 VSS.n498 VSS.n495 5.2005
R2040 VSS.n767 VSS.n498 5.2005
R2041 VSS.n765 VSS.n764 5.2005
R2042 VSS.n766 VSS.n765 5.2005
R2043 VSS.n763 VSS.n505 5.2005
R2044 VSS.n509 VSS.n505 5.2005
R2045 VSS.n762 VSS.n761 5.2005
R2046 VSS.n761 VSS.n760 5.2005
R2047 VSS.n507 VSS.n506 5.2005
R2048 VSS.n752 VSS.n507 5.2005
R2049 VSS.n750 VSS.n749 5.2005
R2050 VSS.n751 VSS.n750 5.2005
R2051 VSS.n748 VSS.n514 5.2005
R2052 VSS.n743 VSS.n514 5.2005
R2053 VSS.n747 VSS.n746 5.2005
R2054 VSS.n746 VSS.n745 5.2005
R2055 VSS.n516 VSS.n515 5.2005
R2056 VSS.n517 VSS.n516 5.2005
R2057 VSS.n552 VSS.n551 5.2005
R2058 VSS.n551 VSS.n550 5.2005
R2059 VSS.n554 VSS.n553 5.2005
R2060 VSS.n556 VSS.n548 5.2005
R2061 VSS.n558 VSS.n557 5.2005
R2062 VSS.n559 VSS.n547 5.2005
R2063 VSS.n561 VSS.n560 5.2005
R2064 VSS.n563 VSS.n546 5.2005
R2065 VSS.n564 VSS.n544 5.2005
R2066 VSS.n567 VSS.n566 5.2005
R2067 VSS.n1810 VSS.n1809 5.2005
R2068 VSS.n1809 VSS.n1808 5.2005
R2069 VSS.n213 VSS.n212 5.2005
R2070 VSS.n1807 VSS.n213 5.2005
R2071 VSS.n1805 VSS.n1804 5.2005
R2072 VSS.n1806 VSS.n1805 5.2005
R2073 VSS.n1803 VSS.n215 5.2005
R2074 VSS.n215 VSS.n214 5.2005
R2075 VSS.n1802 VSS.n1801 5.2005
R2076 VSS.n1801 VSS.n1800 5.2005
R2077 VSS.n217 VSS.n216 5.2005
R2078 VSS.n1799 VSS.n217 5.2005
R2079 VSS.n1797 VSS.n1796 5.2005
R2080 VSS.n1798 VSS.n1797 5.2005
R2081 VSS.n1795 VSS.n219 5.2005
R2082 VSS.n219 VSS.n218 5.2005
R2083 VSS.n1794 VSS.n1793 5.2005
R2084 VSS.n1793 VSS.n1792 5.2005
R2085 VSS.n221 VSS.n220 5.2005
R2086 VSS.n1791 VSS.n221 5.2005
R2087 VSS.n1788 VSS.n1787 5.2005
R2088 VSS.n1789 VSS.n1788 5.2005
R2089 VSS.n1786 VSS.n226 5.2005
R2090 VSS.n226 VSS.n225 5.2005
R2091 VSS.n1785 VSS.n1784 5.2005
R2092 VSS.n1784 VSS.n1783 5.2005
R2093 VSS.n228 VSS.n227 5.2005
R2094 VSS.n1782 VSS.n228 5.2005
R2095 VSS.n1780 VSS.n1779 5.2005
R2096 VSS.n1781 VSS.n1780 5.2005
R2097 VSS.n1778 VSS.n230 5.2005
R2098 VSS.n230 VSS.n229 5.2005
R2099 VSS.n1777 VSS.n1776 5.2005
R2100 VSS.n1776 VSS.n1775 5.2005
R2101 VSS.n2015 VSS.n139 5.2005
R2102 VSS.n145 VSS.n139 5.2005
R2103 VSS.n2017 VSS.n2016 5.2005
R2104 VSS.n2018 VSS.n2017 5.2005
R2105 VSS.n137 VSS.n136 5.2005
R2106 VSS.n2019 VSS.n137 5.2005
R2107 VSS.n2022 VSS.n2021 5.2005
R2108 VSS.n2021 VSS.n2020 5.2005
R2109 VSS.n2023 VSS.n134 5.2005
R2110 VSS.n134 VSS.n132 5.2005
R2111 VSS.n2025 VSS.n2024 5.2005
R2112 VSS.n2026 VSS.n2025 5.2005
R2113 VSS.n135 VSS.n133 5.2005
R2114 VSS.n133 VSS.n131 5.2005
R2115 VSS.n1826 VSS.n1825 5.2005
R2116 VSS.n1827 VSS.n1826 5.2005
R2117 VSS.n1824 VSS.n1823 5.2005
R2118 VSS.n1828 VSS.n1824 5.2005
R2119 VSS.n1831 VSS.n1830 5.2005
R2120 VSS.n1830 VSS.n1829 5.2005
R2121 VSS.n1832 VSS.n1822 5.2005
R2122 VSS.n1822 VSS.n1821 5.2005
R2123 VSS.n1834 VSS.n1833 5.2005
R2124 VSS.n1835 VSS.n1834 5.2005
R2125 VSS.n1820 VSS.n1819 5.2005
R2126 VSS.n1836 VSS.n1820 5.2005
R2127 VSS.n1839 VSS.n1838 5.2005
R2128 VSS.n1838 VSS.n1837 5.2005
R2129 VSS.n1840 VSS.n1818 5.2005
R2130 VSS.n1818 VSS.n1817 5.2005
R2131 VSS.n1842 VSS.n1841 5.2005
R2132 VSS.n1843 VSS.n1842 5.2005
R2133 VSS.n1816 VSS.n1815 5.2005
R2134 VSS.n1844 VSS.n1816 5.2005
R2135 VSS.n1847 VSS.n1846 5.2005
R2136 VSS.n1846 VSS.n1845 5.2005
R2137 VSS.n1848 VSS.n1814 5.2005
R2138 VSS.n1814 VSS.n1813 5.2005
R2139 VSS.n1850 VSS.n1849 5.2005
R2140 VSS.n1851 VSS.n1850 5.2005
R2141 VSS.n1812 VSS.n1811 5.2005
R2142 VSS.n1852 VSS.n1812 5.2005
R2143 VSS.n1855 VSS.n1854 5.2005
R2144 VSS.n1854 VSS.n1853 5.2005
R2145 VSS.n2348 VSS.n2347 5.2005
R2146 VSS.n2207 VSS.n23 5.2005
R2147 VSS.n2209 VSS.n2208 5.2005
R2148 VSS.n2210 VSS.n2205 5.2005
R2149 VSS.n2212 VSS.n2211 5.2005
R2150 VSS.n2214 VSS.n2204 5.2005
R2151 VSS.n2215 VSS.n2203 5.2005
R2152 VSS.n2215 VSS.n27 5.2005
R2153 VSS.n2218 VSS.n2217 5.2005
R2154 VSS.n2217 VSS.n2216 5.2005
R2155 VSS.n2219 VSS.n2202 5.2005
R2156 VSS.n2202 VSS.n2201 5.2005
R2157 VSS.n2221 VSS.n2220 5.2005
R2158 VSS.n2222 VSS.n2221 5.2005
R2159 VSS.n2200 VSS.n2199 5.2005
R2160 VSS.n2223 VSS.n2200 5.2005
R2161 VSS.n2226 VSS.n2225 5.2005
R2162 VSS.n2225 VSS.n2224 5.2005
R2163 VSS.n2227 VSS.n82 5.2005
R2164 VSS.n82 VSS.n80 5.2005
R2165 VSS.n2229 VSS.n2228 5.2005
R2166 VSS.n2230 VSS.n2229 5.2005
R2167 VSS.n2198 VSS.n81 5.2005
R2168 VSS.n81 VSS.n79 5.2005
R2169 VSS.n2197 VSS.n2196 5.2005
R2170 VSS.n2196 VSS.n2195 5.2005
R2171 VSS.n84 VSS.n83 5.2005
R2172 VSS.n2194 VSS.n84 5.2005
R2173 VSS.n2192 VSS.n2191 5.2005
R2174 VSS.n2193 VSS.n2192 5.2005
R2175 VSS.n2190 VSS.n86 5.2005
R2176 VSS.n86 VSS.n85 5.2005
R2177 VSS.n2188 VSS.n2187 5.2005
R2178 VSS.n2187 VSS.n2186 5.2005
R2179 VSS.n90 VSS.n89 5.2005
R2180 VSS.n92 VSS.n90 5.2005
R2181 VSS.n2038 VSS.n2037 5.2005
R2182 VSS.n2039 VSS.n2038 5.2005
R2183 VSS.n2042 VSS.n2041 5.2005
R2184 VSS.n2041 VSS.n2040 5.2005
R2185 VSS.n2043 VSS.n2036 5.2005
R2186 VSS.n2036 VSS.n2035 5.2005
R2187 VSS.n2045 VSS.n2044 5.2005
R2188 VSS.n2046 VSS.n2045 5.2005
R2189 VSS.n2034 VSS.n2033 5.2005
R2190 VSS.n2047 VSS.n2034 5.2005
R2191 VSS.n2050 VSS.n2049 5.2005
R2192 VSS.n2049 VSS.n2048 5.2005
R2193 VSS.n2051 VSS.n125 5.2005
R2194 VSS.n125 VSS.n123 5.2005
R2195 VSS.n2053 VSS.n2052 5.2005
R2196 VSS.n2054 VSS.n2053 5.2005
R2197 VSS.n2032 VSS.n124 5.2005
R2198 VSS.n124 VSS.n122 5.2005
R2199 VSS.n2031 VSS.n2030 5.2005
R2200 VSS.n127 VSS.n126 5.2005
R2201 VSS.n1860 VSS.n1859 5.2005
R2202 VSS.n1861 VSS.n1858 5.2005
R2203 VSS.n1863 VSS.n1862 5.2005
R2204 VSS.n1865 VSS.n1857 5.2005
R2205 VSS.n1866 VSS.n1856 5.2005
R2206 VSS.n1869 VSS.n1868 5.2005
R2207 VSS.n1872 VSS.n1871 5.2005
R2208 VSS.n1874 VSS.n209 5.2005
R2209 VSS.n1876 VSS.n1875 5.2005
R2210 VSS.n1877 VSS.n208 5.2005
R2211 VSS.n1879 VSS.n1878 5.2005
R2212 VSS.n1881 VSS.n205 5.2005
R2213 VSS.n1883 VSS.n1882 5.2005
R2214 VSS.n1884 VSS.n203 5.2005
R2215 VSS.n1886 VSS.n1885 5.2005
R2216 VSS.n204 VSS.n202 5.2005
R2217 VSS.n1889 VSS.n200 5.2005
R2218 VSS.n1889 VSS.n1888 5.2005
R2219 VSS.n1891 VSS.n1890 5.2005
R2220 VSS.n1892 VSS.n199 5.2005
R2221 VSS.n1894 VSS.n1893 5.2005
R2222 VSS.n1896 VSS.n197 5.2005
R2223 VSS.n1898 VSS.n1897 5.2005
R2224 VSS.n1899 VSS.n196 5.2005
R2225 VSS.n1901 VSS.n1900 5.2005
R2226 VSS.n1903 VSS.n194 5.2005
R2227 VSS.n1602 VSS.n193 5.2005
R2228 VSS.n1603 VSS.n1601 5.2005
R2229 VSS.n1605 VSS.n1604 5.2005
R2230 VSS.n1607 VSS.n1598 5.2005
R2231 VSS.n1609 VSS.n1608 5.2005
R2232 VSS.n1610 VSS.n1597 5.2005
R2233 VSS.n1612 VSS.n1611 5.2005
R2234 VSS.n1614 VSS.n1596 5.2005
R2235 VSS.n1615 VSS.n1594 5.2005
R2236 VSS.n1618 VSS.n1617 5.2005
R2237 VSS.n1619 VSS.n1593 5.2005
R2238 VSS.n1595 VSS.n1593 5.2005
R2239 VSS.n1621 VSS.n1620 5.2005
R2240 VSS.n1623 VSS.n1591 5.2005
R2241 VSS.n1625 VSS.n1624 5.2005
R2242 VSS.n1626 VSS.n1590 5.2005
R2243 VSS.n1628 VSS.n1627 5.2005
R2244 VSS.n1630 VSS.n1589 5.2005
R2245 VSS.n1631 VSS.n1588 5.2005
R2246 VSS.n1634 VSS.n1633 5.2005
R2247 VSS.n1587 VSS.n1586 5.2005
R2248 VSS.n1584 VSS.n282 5.2005
R2249 VSS.n1583 VSS.n1582 5.2005
R2250 VSS.n1581 VSS.n1580 5.2005
R2251 VSS.n1579 VSS.n284 5.2005
R2252 VSS.n1577 VSS.n1576 5.2005
R2253 VSS.n1575 VSS.n285 5.2005
R2254 VSS.n1574 VSS.n1573 5.2005
R2255 VSS.n1571 VSS.n286 5.2005
R2256 VSS.n1566 VSS.n287 5.2005
R2257 VSS.n1568 VSS.n1567 5.2005
R2258 VSS.n1569 VSS.n1568 5.2005
R2259 VSS.n1565 VSS.n288 5.2005
R2260 VSS.n1564 VSS.n1563 5.2005
R2261 VSS.n290 VSS.n289 5.2005
R2262 VSS.n1559 VSS.n1558 5.2005
R2263 VSS.n1557 VSS.n298 5.2005
R2264 VSS.n1556 VSS.n1555 5.2005
R2265 VSS.n1554 VSS.n1553 5.2005
R2266 VSS.n1552 VSS.n1551 5.2005
R2267 VSS.n1549 VSS.n1548 5.2005
R2268 VSS.n1547 VSS.n1546 5.2005
R2269 VSS.n1545 VSS.n1544 5.2005
R2270 VSS.n1543 VSS.n1542 5.2005
R2271 VSS.n1541 VSS.n1540 5.2005
R2272 VSS.n1539 VSS.n1538 5.2005
R2273 VSS.n1537 VSS.n1536 5.2005
R2274 VSS.n1535 VSS.n1534 5.2005
R2275 VSS.n1533 VSS.n302 5.2005
R2276 VSS.n1528 VSS.n303 5.2005
R2277 VSS.n1530 VSS.n1529 5.2005
R2278 VSS.n1531 VSS.n1530 5.2005
R2279 VSS.n1527 VSS.n304 5.2005
R2280 VSS.n1526 VSS.n1525 5.2005
R2281 VSS.n306 VSS.n305 5.2005
R2282 VSS.n1521 VSS.n1520 5.2005
R2283 VSS.n1519 VSS.n314 5.2005
R2284 VSS.n1518 VSS.n1517 5.2005
R2285 VSS.n1516 VSS.n1515 5.2005
R2286 VSS.n1514 VSS.n1513 5.2005
R2287 VSS.n1511 VSS.n1510 5.2005
R2288 VSS.n1509 VSS.n1508 5.2005
R2289 VSS.n1507 VSS.n1506 5.2005
R2290 VSS.n1505 VSS.n1504 5.2005
R2291 VSS.n1503 VSS.n1502 5.2005
R2292 VSS.n1501 VSS.n1500 5.2005
R2293 VSS.n1499 VSS.n1498 5.2005
R2294 VSS.n1497 VSS.n1496 5.2005
R2295 VSS.n1495 VSS.n318 5.2005
R2296 VSS.n1490 VSS.n319 5.2005
R2297 VSS.n1492 VSS.n1491 5.2005
R2298 VSS.n1493 VSS.n1492 5.2005
R2299 VSS.n1489 VSS.n320 5.2005
R2300 VSS.n324 VSS.n320 5.2005
R2301 VSS.n1488 VSS.n1487 5.2005
R2302 VSS.n1487 VSS.n1486 5.2005
R2303 VSS.n322 VSS.n321 5.2005
R2304 VSS.n1138 VSS.n322 5.2005
R2305 VSS.n1144 VSS.n1143 5.2005
R2306 VSS.n1145 VSS.n1144 5.2005
R2307 VSS.n1142 VSS.n1140 5.2005
R2308 VSS.n1140 VSS.n1137 5.2005
R2309 VSS.n1141 VSS.n822 5.2005
R2310 VSS.n824 VSS.n822 5.2005
R2311 VSS.n1154 VSS.n821 5.2005
R2312 VSS.n1154 VSS.n1153 5.2005
R2313 VSS.n1156 VSS.n1155 5.2005
R2314 VSS.n1155 VSS.n492 5.2005
R2315 VSS.n1159 VSS.n1158 5.2005
R2316 VSS.n1160 VSS.n1159 5.2005
R2317 VSS.n771 VSS.n500 5.2005
R2318 VSS.n500 VSS.n499 5.2005
R2319 VSS.n770 VSS.n769 5.2005
R2320 VSS.n769 VSS.n768 5.2005
R2321 VSS.n503 VSS.n502 5.2005
R2322 VSS.n504 VSS.n503 5.2005
R2323 VSS.n758 VSS.n757 5.2005
R2324 VSS.n759 VSS.n758 5.2005
R2325 VSS.n756 VSS.n510 5.2005
R2326 VSS.n510 VSS.n508 5.2005
R2327 VSS.n755 VSS.n754 5.2005
R2328 VSS.n754 VSS.n753 5.2005
R2329 VSS.n512 VSS.n511 5.2005
R2330 VSS.n742 VSS.n512 5.2005
R2331 VSS.n612 VSS.n611 5.2005
R2332 VSS.n614 VSS.n610 5.2005
R2333 VSS.n615 VSS.n608 5.2005
R2334 VSS.n615 VSS.n521 5.2005
R2335 VSS.n617 VSS.n616 5.2005
R2336 VSS.n618 VSS.n607 5.2005
R2337 VSS.n620 VSS.n619 5.2005
R2338 VSS.n622 VSS.n605 5.2005
R2339 VSS.n624 VSS.n623 5.2005
R2340 VSS.n625 VSS.n604 5.2005
R2341 VSS.n627 VSS.n626 5.2005
R2342 VSS.n629 VSS.n603 5.2005
R2343 VSS.n48 VSS.n47 5.2005
R2344 VSS.n2303 VSS.n48 5.2005
R2345 VSS.n2306 VSS.n2305 5.2005
R2346 VSS.n2305 VSS.n2304 5.2005
R2347 VSS.n2307 VSS.n46 5.2005
R2348 VSS.n46 VSS.n45 5.2005
R2349 VSS.n2309 VSS.n2308 5.2005
R2350 VSS.n2310 VSS.n2309 5.2005
R2351 VSS.n44 VSS.n43 5.2005
R2352 VSS.n2311 VSS.n44 5.2005
R2353 VSS.n2314 VSS.n2313 5.2005
R2354 VSS.n2313 VSS.n2312 5.2005
R2355 VSS.n2315 VSS.n42 5.2005
R2356 VSS.n42 VSS.n41 5.2005
R2357 VSS.n2317 VSS.n2316 5.2005
R2358 VSS.n2318 VSS.n2317 5.2005
R2359 VSS.n40 VSS.n39 5.2005
R2360 VSS.n2319 VSS.n40 5.2005
R2361 VSS.n2322 VSS.n2321 5.2005
R2362 VSS.n2321 VSS.n2320 5.2005
R2363 VSS.n2323 VSS.n38 5.2005
R2364 VSS.n38 VSS.n37 5.2005
R2365 VSS.n2325 VSS.n2324 5.2005
R2366 VSS.n2326 VSS.n2325 5.2005
R2367 VSS.n36 VSS.n35 5.2005
R2368 VSS.n2327 VSS.n36 5.2005
R2369 VSS.n2330 VSS.n2329 5.2005
R2370 VSS.n2329 VSS.n2328 5.2005
R2371 VSS.n2331 VSS.n34 5.2005
R2372 VSS.n34 VSS.n33 5.2005
R2373 VSS.n2333 VSS.n2332 5.2005
R2374 VSS.n2334 VSS.n2333 5.2005
R2375 VSS.n32 VSS.n31 5.2005
R2376 VSS.n2335 VSS.n32 5.2005
R2377 VSS.n2338 VSS.n2337 5.2005
R2378 VSS.n2337 VSS.n2336 5.2005
R2379 VSS.n2339 VSS.n29 5.2005
R2380 VSS.n29 VSS.n28 5.2005
R2381 VSS.n2341 VSS.n2340 5.2005
R2382 VSS.n2342 VSS.n2341 5.2005
R2383 VSS.n30 VSS.n25 5.2005
R2384 VSS.n2343 VSS.n25 5.2005
R2385 VSS.n2345 VSS.n22 5.2005
R2386 VSS.n2345 VSS.n2344 5.2005
R2387 VSS.n2299 VSS.n2298 5.2005
R2388 VSS.n52 VSS.n51 5.2005
R2389 VSS.n2249 VSS.n2248 5.2005
R2390 VSS.n2250 VSS.n2247 5.2005
R2391 VSS.n2252 VSS.n2251 5.2005
R2392 VSS.n2252 VSS.n49 5.2005
R2393 VSS.n2253 VSS.n2246 5.2005
R2394 VSS.n2254 VSS.n2253 5.2005
R2395 VSS.n2257 VSS.n2256 5.2005
R2396 VSS.n2256 VSS.n2255 5.2005
R2397 VSS.n2258 VSS.n2245 5.2005
R2398 VSS.n2245 VSS.n2244 5.2005
R2399 VSS.n2260 VSS.n2259 5.2005
R2400 VSS.n2261 VSS.n2260 5.2005
R2401 VSS.n2243 VSS.n2242 5.2005
R2402 VSS.n2262 VSS.n2243 5.2005
R2403 VSS.n2265 VSS.n2264 5.2005
R2404 VSS.n2264 VSS.n2263 5.2005
R2405 VSS.n2266 VSS.n2234 5.2005
R2406 VSS.n2234 VSS.n2233 5.2005
R2407 VSS.n2268 VSS.n2267 5.2005
R2408 VSS.n2269 VSS.n2268 5.2005
R2409 VSS.n2241 VSS.n2232 5.2005
R2410 VSS.n2240 VSS.n2239 5.2005
R2411 VSS.n2238 VSS.n2237 5.2005
R2412 VSS.n2236 VSS.n2235 5.2005
R2413 VSS.n62 VSS.n55 5.2005
R2414 VSS.n58 VSS.n54 5.2005
R2415 VSS.n2288 VSS.n2287 5.2005
R2416 VSS.n2290 VSS.n2289 5.2005
R2417 VSS.n2291 VSS.n67 5.2005
R2418 VSS.n2293 VSS.n2292 5.2005
R2419 VSS.n2294 VSS.n2293 5.2005
R2420 VSS.n2286 VSS.n66 5.2005
R2421 VSS.n2282 VSS.n66 5.2005
R2422 VSS.n2285 VSS.n2284 5.2005
R2423 VSS.n2284 VSS.n2283 5.2005
R2424 VSS.n69 VSS.n68 5.2005
R2425 VSS.n70 VSS.n69 5.2005
R2426 VSS.n1997 VSS.n1994 5.2005
R2427 VSS.n1994 VSS.n1993 5.2005
R2428 VSS.n1999 VSS.n1998 5.2005
R2429 VSS.n2000 VSS.n1999 5.2005
R2430 VSS.n1995 VSS.n1992 5.2005
R2431 VSS.n2001 VSS.n1992 5.2005
R2432 VSS.n2003 VSS.n1990 5.2005
R2433 VSS.n2003 VSS.n2002 5.2005
R2434 VSS.n2005 VSS.n2004 5.2005
R2435 VSS.n2006 VSS.n1988 5.2005
R2436 VSS.n2008 VSS.n2007 5.2005
R2437 VSS.n1989 VSS.n1987 5.2005
R2438 VSS.n1986 VSS.n141 5.2005
R2439 VSS.n2014 VSS.n142 5.2005
R2440 VSS.n2014 VSS.n2013 5.2005
R2441 VSS.n144 VSS.n140 5.2005
R2442 VSS.n1983 VSS.n1982 5.2005
R2443 VSS.n1981 VSS.n147 5.2005
R2444 VSS.n1980 VSS.n1979 5.2005
R2445 VSS.n1978 VSS.n1977 5.2005
R2446 VSS.n1976 VSS.n148 5.2005
R2447 VSS.n1976 VSS.n1975 5.2005
R2448 VSS.n1970 VSS.n149 5.2005
R2449 VSS.n1974 VSS.n149 5.2005
R2450 VSS.n1972 VSS.n1971 5.2005
R2451 VSS.n1973 VSS.n1972 5.2005
R2452 VSS.n1969 VSS.n151 5.2005
R2453 VSS.n151 VSS.n150 5.2005
R2454 VSS.n1968 VSS.n1967 5.2005
R2455 VSS.n1967 VSS.n1966 5.2005
R2456 VSS.n155 VSS.n152 5.2005
R2457 VSS.n1965 VSS.n155 5.2005
R2458 VSS.n1963 VSS.n1962 5.2005
R2459 VSS.n1964 VSS.n1963 5.2005
R2460 VSS.n1961 VSS.n157 5.2005
R2461 VSS.n1960 VSS.n1959 5.2005
R2462 VSS.n159 VSS.n158 5.2005
R2463 VSS.n1955 VSS.n1954 5.2005
R2464 VSS.n1953 VSS.n165 5.2005
R2465 VSS.n1952 VSS.n168 5.2005
R2466 VSS.n1952 VSS.n1951 5.2005
R2467 VSS.n1413 VSS.n166 5.2005
R2468 VSS.n1415 VSS.n1414 5.2005
R2469 VSS.n1417 VSS.n1416 5.2005
R2470 VSS.n1419 VSS.n1418 5.2005
R2471 VSS.n1421 VSS.n1420 5.2005
R2472 VSS.n1422 VSS.n1412 5.2005
R2473 VSS.n1423 VSS.n1422 5.2005
R2474 VSS.n1426 VSS.n1425 5.2005
R2475 VSS.n1425 VSS.n1424 5.2005
R2476 VSS.n1427 VSS.n1411 5.2005
R2477 VSS.n1411 VSS.n1410 5.2005
R2478 VSS.n1429 VSS.n1428 5.2005
R2479 VSS.n1430 VSS.n1429 5.2005
R2480 VSS.n1408 VSS.n1407 5.2005
R2481 VSS.n1431 VSS.n1408 5.2005
R2482 VSS.n1434 VSS.n1433 5.2005
R2483 VSS.n1433 VSS.n1432 5.2005
R2484 VSS.n1435 VSS.n367 5.2005
R2485 VSS.n1409 VSS.n367 5.2005
R2486 VSS.n1437 VSS.n1436 5.2005
R2487 VSS.n374 VSS.n366 5.2005
R2488 VSS.n373 VSS.n372 5.2005
R2489 VSS.n371 VSS.n370 5.2005
R2490 VSS.n369 VSS.n368 5.2005
R2491 VSS.n363 VSS.n356 5.2005
R2492 VSS.n361 VSS.n356 5.2005
R2493 VSS.n1282 VSS.n1281 5.2005
R2494 VSS.n1284 VSS.n1283 5.2005
R2495 VSS.n1286 VSS.n1285 5.2005
R2496 VSS.n1288 VSS.n1287 5.2005
R2497 VSS.n1290 VSS.n1289 5.2005
R2498 VSS.n1291 VSS.n1280 5.2005
R2499 VSS.n1292 VSS.n1291 5.2005
R2500 VSS.n1295 VSS.n1294 5.2005
R2501 VSS.n1294 VSS.n1293 5.2005
R2502 VSS.n1296 VSS.n1279 5.2005
R2503 VSS.n1279 VSS.n1278 5.2005
R2504 VSS.n1298 VSS.n1297 5.2005
R2505 VSS.n1299 VSS.n1298 5.2005
R2506 VSS.n1277 VSS.n377 5.2005
R2507 VSS.n1300 VSS.n1277 5.2005
R2508 VSS.n1303 VSS.n1302 5.2005
R2509 VSS.n1302 VSS.n1301 5.2005
R2510 VSS.n1304 VSS.n1276 5.2005
R2511 VSS.n1276 VSS.n1255 5.2005
R2512 VSS.n1306 VSS.n1305 5.2005
R2513 VSS.n1308 VSS.n1274 5.2005
R2514 VSS.n1310 VSS.n1309 5.2005
R2515 VSS.n1311 VSS.n1273 5.2005
R2516 VSS.n1313 VSS.n1312 5.2005
R2517 VSS.n1315 VSS.n378 5.2005
R2518 VSS.n1272 VSS.n378 5.2005
R2519 VSS.n1270 VSS.n1269 5.2005
R2520 VSS.n1268 VSS.n1259 5.2005
R2521 VSS.n1267 VSS.n1266 5.2005
R2522 VSS.n1264 VSS.n1260 5.2005
R2523 VSS.n1262 VSS.n1261 5.2005
R2524 VSS.n1254 VSS.n1253 5.2005
R2525 VSS.n1379 VSS.n1254 5.2005
R2526 VSS.n1382 VSS.n1381 5.2005
R2527 VSS.n1381 VSS.n1380 5.2005
R2528 VSS.n1383 VSS.n1252 5.2005
R2529 VSS.n1252 VSS.n1251 5.2005
R2530 VSS.n1385 VSS.n1384 5.2005
R2531 VSS.n1386 VSS.n1385 5.2005
R2532 VSS.n1249 VSS.n380 5.2005
R2533 VSS.n1387 VSS.n1249 5.2005
R2534 VSS.n1390 VSS.n1389 5.2005
R2535 VSS.n1389 VSS.n1388 5.2005
R2536 VSS.n1391 VSS.n1242 5.2005
R2537 VSS.n1250 VSS.n1242 5.2005
R2538 VSS.n1393 VSS.n1392 5.2005
R2539 VSS.n1248 VSS.n1241 5.2005
R2540 VSS.n1247 VSS.n1246 5.2005
R2541 VSS.n1245 VSS.n1244 5.2005
R2542 VSS.n1243 VSS.n383 5.2005
R2543 VSS.n1400 VSS.n385 5.2005
R2544 VSS.n1400 VSS.n1399 5.2005
R2545 VSS.n450 VSS.n382 5.2005
R2546 VSS.n1237 VSS.n1236 5.2005
R2547 VSS.n1235 VSS.n449 5.2005
R2548 VSS.n1234 VSS.n1233 5.2005
R2549 VSS.n1232 VSS.n1231 5.2005
R2550 VSS.n1230 VSS.n451 5.2005
R2551 VSS.n1230 VSS.n1229 5.2005
R2552 VSS.n1224 VSS.n452 5.2005
R2553 VSS.n1228 VSS.n452 5.2005
R2554 VSS.n1226 VSS.n1225 5.2005
R2555 VSS.n1227 VSS.n1226 5.2005
R2556 VSS.n1223 VSS.n454 5.2005
R2557 VSS.n454 VSS.n453 5.2005
R2558 VSS.n1222 VSS.n1221 5.2005
R2559 VSS.n1221 VSS.n1220 5.2005
R2560 VSS.n457 VSS.n455 5.2005
R2561 VSS.n1219 VSS.n457 5.2005
R2562 VSS.n1217 VSS.n1216 5.2005
R2563 VSS.n1218 VSS.n1217 5.2005
R2564 VSS.n1215 VSS.n459 5.2005
R2565 VSS.n1214 VSS.n1213 5.2005
R2566 VSS.n461 VSS.n460 5.2005
R2567 VSS.n1209 VSS.n1208 5.2005
R2568 VSS.n1207 VSS.n467 5.2005
R2569 VSS.n1206 VSS.n470 5.2005
R2570 VSS.n1206 VSS.n1205 5.2005
R2571 VSS.n674 VSS.n468 5.2005
R2572 VSS.n676 VSS.n675 5.2005
R2573 VSS.n678 VSS.n677 5.2005
R2574 VSS.n680 VSS.n679 5.2005
R2575 VSS.n682 VSS.n681 5.2005
R2576 VSS.n683 VSS.n673 5.2005
R2577 VSS.n684 VSS.n683 5.2005
R2578 VSS.n687 VSS.n686 5.2005
R2579 VSS.n686 VSS.n685 5.2005
R2580 VSS.n688 VSS.n672 5.2005
R2581 VSS.n672 VSS.n671 5.2005
R2582 VSS.n690 VSS.n689 5.2005
R2583 VSS.n691 VSS.n690 5.2005
R2584 VSS.n669 VSS.n668 5.2005
R2585 VSS.n692 VSS.n669 5.2005
R2586 VSS.n695 VSS.n694 5.2005
R2587 VSS.n694 VSS.n693 5.2005
R2588 VSS.n696 VSS.n658 5.2005
R2589 VSS.n670 VSS.n658 5.2005
R2590 VSS.n698 VSS.n697 5.2005
R2591 VSS.n665 VSS.n657 5.2005
R2592 VSS.n664 VSS.n663 5.2005
R2593 VSS.n662 VSS.n661 5.2005
R2594 VSS.n660 VSS.n659 5.2005
R2595 VSS.n653 VSS.n652 5.2005
R2596 VSS.n2173 VSS.n2164 5.2005
R2597 VSS.n2164 VSS.n2163 5.2005
R2598 VSS.n2175 VSS.n2174 5.2005
R2599 VSS.n2176 VSS.n2175 5.2005
R2600 VSS.n2162 VSS.n2161 5.2005
R2601 VSS.n2177 VSS.n2162 5.2005
R2602 VSS.n2180 VSS.n2179 5.2005
R2603 VSS.n2179 VSS.n2178 5.2005
R2604 VSS.n2181 VSS.n2142 5.2005
R2605 VSS.n2142 VSS.n2140 5.2005
R2606 VSS.n2183 VSS.n2182 5.2005
R2607 VSS.n2184 VSS.n2183 5.2005
R2608 VSS.n2160 VSS.n2141 5.2005
R2609 VSS.n2159 VSS.n2158 5.2005
R2610 VSS.n2156 VSS.n2143 5.2005
R2611 VSS.n2154 VSS.n2153 5.2005
R2612 VSS.n2152 VSS.n2144 5.2005
R2613 VSS.n2151 VSS.n2150 5.2005
R2614 VSS.n2148 VSS.n2145 5.2005
R2615 VSS.n2146 VSS.n87 5.2005
R2616 VSS.n2172 VSS.n2166 5.2005
R2617 VSS.n2166 VSS.n2165 5.2005
R2618 VSS.n74 VSS.n56 5.2005
R2619 VSS.n74 VSS.n60 5.2005
R2620 VSS.n2277 VSS.n75 5.2005
R2621 VSS.n75 VSS.n72 5.2005
R2622 VSS.n2279 VSS.n2278 5.2005
R2623 VSS.n2280 VSS.n2279 5.2005
R2624 VSS.n2276 VSS.n73 5.2005
R2625 VSS.n73 VSS.n71 5.2005
R2626 VSS.n2275 VSS.n2274 5.2005
R2627 VSS.n2274 VSS.n2273 5.2005
R2628 VSS.n77 VSS.n76 5.2005
R2629 VSS.n2272 VSS.n77 5.2005
R2630 VSS.n2171 VSS.n2170 5.2005
R2631 VSS.n2170 VSS.n78 5.2005
R2632 VSS.n2296 VSS.n57 5.2005
R2633 VSS.n2294 VSS.n57 5.2005
R2634 VSS.n2296 VSS.n2295 5.2005
R2635 VSS.n2295 VSS.n2294 5.2005
R2636 VSS.n2384 VSS.n2 5.06478
R2637 VSS.n1167 VSS.n490 4.93804
R2638 VSS.n2169 VSS.n2167 4.55948
R2639 VSS.n2169 VSS.n2168 4.38259
R2640 VSS.n740 VSS.n522 4.18325
R2641 VSS.n1479 VSS.n330 4.05793
R2642 VSS.n1481 VSS.n328 4.05793
R2643 VSS.n1483 VSS.n326 4.05793
R2644 VSS.n1168 VSS.n1167 4.05793
R2645 VSS.n1914 VSS.n1913 4.05793
R2646 VSS.n2346 VSS.n21 3.59261
R2647 VSS.n96 VSS.n91 3.59261
R2648 VSS.n1904 VSS.n192 3.59261
R2649 VSS.n1637 VSS.n280 3.59261
R2650 VSS.n1550 VSS.n300 3.59261
R2651 VSS.n1512 VSS.n316 3.59261
R2652 VSS.n811 VSS.n501 3.59261
R2653 VSS.n630 VSS.n527 3.59261
R2654 VSS.n1809 VSS.n211 3.59261
R2655 VSS.n2378 VSS.n4 3.32459
R2656 VSS.n2374 VSS.n3 3.32459
R2657 VSS.n2132 VSS.n93 3.32459
R2658 VSS.n2128 VSS.n94 3.32459
R2659 VSS.n2124 VSS.n95 3.32459
R2660 VSS.n97 VSS.n96 3.32459
R2661 VSS.n781 VSS.n779 3.32459
R2662 VSS.n788 VSS.n787 3.32459
R2663 VSS.n789 VSS.n777 3.32459
R2664 VSS.n796 VSS.n795 3.32459
R2665 VSS.n797 VSS.n775 3.32459
R2666 VSS.n804 VSS.n803 3.32459
R2667 VSS.n808 VSS.n773 3.32459
R2668 VSS.n811 VSS.n810 3.32459
R2669 VSS.n819 VSS.n818 3.32459
R2670 VSS.n816 VSS.n814 3.32459
R2671 VSS.n810 VSS.n809 3.32459
R2672 VSS.n805 VSS.n773 3.32459
R2673 VSS.n803 VSS.n802 3.32459
R2674 VSS.n798 VSS.n797 3.32459
R2675 VSS.n795 VSS.n794 3.32459
R2676 VSS.n790 VSS.n789 3.32459
R2677 VSS.n787 VSS.n786 3.32459
R2678 VSS.n782 VSS.n781 3.32459
R2679 VSS.n814 VSS.n489 3.32459
R2680 VSS.n818 VSS.n817 3.32459
R2681 VSS.n2123 VSS.n97 3.32459
R2682 VSS.n2127 VSS.n95 3.32459
R2683 VSS.n2131 VSS.n94 3.32459
R2684 VSS.n100 VSS.n93 3.32459
R2685 VSS.n2377 VSS.n3 3.32459
R2686 VSS.n6 VSS.n4 3.32459
R2687 VSS.n565 VSS.n564 3.32459
R2688 VSS.n562 VSS.n561 3.32459
R2689 VSS.n557 VSS.n549 3.32459
R2690 VSS.n555 VSS.n554 3.32459
R2691 VSS.n1128 VSS.n1127 3.32459
R2692 VSS.n1123 VSS.n832 3.32459
R2693 VSS.n1121 VSS.n1120 3.32459
R2694 VSS.n1116 VSS.n836 3.32459
R2695 VSS.n1114 VSS.n1113 3.32459
R2696 VSS.n1108 VSS.n1107 3.32459
R2697 VSS.n1103 VSS.n892 3.32459
R2698 VSS.n1101 VSS.n1100 3.32459
R2699 VSS.n1096 VSS.n895 3.32459
R2700 VSS.n1093 VSS.n1092 3.32459
R2701 VSS.n1088 VSS.n900 3.32459
R2702 VSS.n1086 VSS.n1085 3.32459
R2703 VSS.n1081 VSS.n904 3.32459
R2704 VSS.n1079 VSS.n1078 3.32459
R2705 VSS.n1073 VSS.n1072 3.32459
R2706 VSS.n1068 VSS.n959 3.32459
R2707 VSS.n1066 VSS.n1065 3.32459
R2708 VSS.n1061 VSS.n962 3.32459
R2709 VSS.n1058 VSS.n1057 3.32459
R2710 VSS.n1053 VSS.n967 3.32459
R2711 VSS.n1051 VSS.n1050 3.32459
R2712 VSS.n1046 VSS.n971 3.32459
R2713 VSS.n1044 VSS.n1043 3.32459
R2714 VSS.n1038 VSS.n1037 3.32459
R2715 VSS.n1033 VSS.n998 3.32459
R2716 VSS.n1031 VSS.n1030 3.32459
R2717 VSS.n1026 VSS.n1001 3.32459
R2718 VSS.n1023 VSS.n1022 3.32459
R2719 VSS.n1018 VSS.n242 3.32459
R2720 VSS.n1014 VSS.n243 3.32459
R2721 VSS.n1010 VSS.n244 3.32459
R2722 VSS.n1005 VSS.n245 3.32459
R2723 VSS.n248 VSS.n246 3.32459
R2724 VSS.n254 VSS.n253 3.32459
R2725 VSS.n1701 VSS.n1700 3.32459
R2726 VSS.n1705 VSS.n239 3.32459
R2727 VSS.n1708 VSS.n237 3.32459
R2728 VSS.n1715 VSS.n1714 3.32459
R2729 VSS.n1716 VSS.n235 3.32459
R2730 VSS.n1723 VSS.n1722 3.32459
R2731 VSS.n1728 VSS.n232 3.32459
R2732 VSS.n1772 VSS.n1771 3.32459
R2733 VSS.n1767 VSS.n1765 3.32459
R2734 VSS.n1762 VSS.n119 3.32459
R2735 VSS.n1758 VSS.n120 3.32459
R2736 VSS.n1754 VSS.n121 3.32459
R2737 VSS.n1751 VSS.n1750 3.32459
R2738 VSS.n1746 VSS.n1736 3.32459
R2739 VSS.n1744 VSS.n1743 3.32459
R2740 VSS.n1738 VSS.n1737 3.32459
R2741 VSS.n2101 VSS.n2100 3.32459
R2742 VSS.n2096 VSS.n114 3.32459
R2743 VSS.n114 VSS.n112 3.32459
R2744 VSS.n2102 VSS.n2101 3.32459
R2745 VSS.n1739 VSS.n1738 3.32459
R2746 VSS.n1745 VSS.n1744 3.32459
R2747 VSS.n1736 VSS.n1734 3.32459
R2748 VSS.n1752 VSS.n1751 3.32459
R2749 VSS.n1757 VSS.n121 3.32459
R2750 VSS.n1761 VSS.n120 3.32459
R2751 VSS.n1766 VSS.n119 3.32459
R2752 VSS.n1765 VSS.n1730 3.32459
R2753 VSS.n1773 VSS.n1772 3.32459
R2754 VSS.n1724 VSS.n232 3.32459
R2755 VSS.n1722 VSS.n1721 3.32459
R2756 VSS.n1717 VSS.n1716 3.32459
R2757 VSS.n1714 VSS.n1713 3.32459
R2758 VSS.n1709 VSS.n1708 3.32459
R2759 VSS.n1702 VSS.n239 3.32459
R2760 VSS.n1700 VSS.n241 3.32459
R2761 VSS.n254 VSS.n247 3.32459
R2762 VSS.n258 VSS.n246 3.32459
R2763 VSS.n1009 VSS.n245 3.32459
R2764 VSS.n1013 VSS.n244 3.32459
R2765 VSS.n1017 VSS.n243 3.32459
R2766 VSS.n1003 VSS.n242 3.32459
R2767 VSS.n1023 VSS.n1002 3.32459
R2768 VSS.n1001 VSS.n999 3.32459
R2769 VSS.n1032 VSS.n1031 3.32459
R2770 VSS.n998 VSS.n996 3.32459
R2771 VSS.n1039 VSS.n1038 3.32459
R2772 VSS.n1045 VSS.n1044 3.32459
R2773 VSS.n971 VSS.n969 3.32459
R2774 VSS.n1052 VSS.n1051 3.32459
R2775 VSS.n967 VSS.n964 3.32459
R2776 VSS.n1058 VSS.n963 3.32459
R2777 VSS.n962 VSS.n960 3.32459
R2778 VSS.n1067 VSS.n1066 3.32459
R2779 VSS.n959 VSS.n957 3.32459
R2780 VSS.n1074 VSS.n1073 3.32459
R2781 VSS.n1080 VSS.n1079 3.32459
R2782 VSS.n904 VSS.n902 3.32459
R2783 VSS.n1087 VSS.n1086 3.32459
R2784 VSS.n900 VSS.n897 3.32459
R2785 VSS.n1093 VSS.n896 3.32459
R2786 VSS.n895 VSS.n893 3.32459
R2787 VSS.n1102 VSS.n1101 3.32459
R2788 VSS.n892 VSS.n890 3.32459
R2789 VSS.n1109 VSS.n1108 3.32459
R2790 VSS.n1115 VSS.n1114 3.32459
R2791 VSS.n836 VSS.n834 3.32459
R2792 VSS.n1122 VSS.n1121 3.32459
R2793 VSS.n832 VSS.n830 3.32459
R2794 VSS.n1128 VSS.n829 3.32459
R2795 VSS.n556 VSS.n555 3.32459
R2796 VSS.n549 VSS.n547 3.32459
R2797 VSS.n563 VSS.n562 3.32459
R2798 VSS.n566 VSS.n565 3.32459
R2799 VSS.n628 VSS.n627 3.32459
R2800 VSS.n623 VSS.n606 3.32459
R2801 VSS.n621 VSS.n620 3.32459
R2802 VSS.n616 VSS.n609 3.32459
R2803 VSS.n613 VSS.n612 3.32459
R2804 VSS.n1495 VSS.n1494 3.32459
R2805 VSS.n1499 VSS.n308 3.32459
R2806 VSS.n1503 VSS.n309 3.32459
R2807 VSS.n1507 VSS.n310 3.32459
R2808 VSS.n1511 VSS.n311 3.32459
R2809 VSS.n1516 VSS.n312 3.32459
R2810 VSS.n314 VSS.n313 3.32459
R2811 VSS.n1522 VSS.n306 3.32459
R2812 VSS.n1524 VSS.n304 3.32459
R2813 VSS.n1533 VSS.n1532 3.32459
R2814 VSS.n1537 VSS.n292 3.32459
R2815 VSS.n1541 VSS.n293 3.32459
R2816 VSS.n1545 VSS.n294 3.32459
R2817 VSS.n1549 VSS.n295 3.32459
R2818 VSS.n1554 VSS.n296 3.32459
R2819 VSS.n298 VSS.n297 3.32459
R2820 VSS.n1560 VSS.n290 3.32459
R2821 VSS.n1562 VSS.n288 3.32459
R2822 VSS.n1571 VSS.n1570 3.32459
R2823 VSS.n1572 VSS.n285 3.32459
R2824 VSS.n1579 VSS.n1578 3.32459
R2825 VSS.n1583 VSS.n283 3.32459
R2826 VSS.n1586 VSS.n1585 3.32459
R2827 VSS.n1632 VSS.n1631 3.32459
R2828 VSS.n1629 VSS.n1628 3.32459
R2829 VSS.n1624 VSS.n1592 3.32459
R2830 VSS.n1622 VSS.n1621 3.32459
R2831 VSS.n1616 VSS.n1615 3.32459
R2832 VSS.n1613 VSS.n1612 3.32459
R2833 VSS.n1608 VSS.n1599 3.32459
R2834 VSS.n1606 VSS.n1605 3.32459
R2835 VSS.n1600 VSS.n193 3.32459
R2836 VSS.n1902 VSS.n1901 3.32459
R2837 VSS.n1897 VSS.n198 3.32459
R2838 VSS.n1895 VSS.n1894 3.32459
R2839 VSS.n1890 VSS.n201 3.32459
R2840 VSS.n1887 VSS.n1886 3.32459
R2841 VSS.n1882 VSS.n206 3.32459
R2842 VSS.n1880 VSS.n1879 3.32459
R2843 VSS.n1875 VSS.n210 3.32459
R2844 VSS.n1873 VSS.n1872 3.32459
R2845 VSS.n1867 VSS.n1866 3.32459
R2846 VSS.n1864 VSS.n1863 3.32459
R2847 VSS.n1859 VSS.n129 3.32459
R2848 VSS.n2030 VSS.n2029 3.32459
R2849 VSS.n2213 VSS.n2212 3.32459
R2850 VSS.n2208 VSS.n2206 3.32459
R2851 VSS.n2347 VSS.n24 3.32459
R2852 VSS.n2207 VSS.n24 3.32459
R2853 VSS.n2206 VSS.n2205 3.32459
R2854 VSS.n2214 VSS.n2213 3.32459
R2855 VSS.n2029 VSS.n127 3.32459
R2856 VSS.n1858 VSS.n129 3.32459
R2857 VSS.n1865 VSS.n1864 3.32459
R2858 VSS.n1868 VSS.n1867 3.32459
R2859 VSS.n1874 VSS.n1873 3.32459
R2860 VSS.n210 VSS.n208 3.32459
R2861 VSS.n1881 VSS.n1880 3.32459
R2862 VSS.n206 VSS.n203 3.32459
R2863 VSS.n1887 VSS.n202 3.32459
R2864 VSS.n201 VSS.n199 3.32459
R2865 VSS.n1896 VSS.n1895 3.32459
R2866 VSS.n198 VSS.n196 3.32459
R2867 VSS.n1903 VSS.n1902 3.32459
R2868 VSS.n1601 VSS.n1600 3.32459
R2869 VSS.n1607 VSS.n1606 3.32459
R2870 VSS.n1599 VSS.n1597 3.32459
R2871 VSS.n1614 VSS.n1613 3.32459
R2872 VSS.n1617 VSS.n1616 3.32459
R2873 VSS.n1623 VSS.n1622 3.32459
R2874 VSS.n1592 VSS.n1590 3.32459
R2875 VSS.n1630 VSS.n1629 3.32459
R2876 VSS.n1633 VSS.n1632 3.32459
R2877 VSS.n1585 VSS.n1584 3.32459
R2878 VSS.n1580 VSS.n283 3.32459
R2879 VSS.n1578 VSS.n1577 3.32459
R2880 VSS.n1573 VSS.n1572 3.32459
R2881 VSS.n1570 VSS.n287 3.32459
R2882 VSS.n1563 VSS.n1562 3.32459
R2883 VSS.n1560 VSS.n1559 3.32459
R2884 VSS.n1555 VSS.n297 3.32459
R2885 VSS.n1551 VSS.n296 3.32459
R2886 VSS.n1546 VSS.n295 3.32459
R2887 VSS.n1542 VSS.n294 3.32459
R2888 VSS.n1538 VSS.n293 3.32459
R2889 VSS.n1534 VSS.n292 3.32459
R2890 VSS.n1532 VSS.n303 3.32459
R2891 VSS.n1525 VSS.n1524 3.32459
R2892 VSS.n1522 VSS.n1521 3.32459
R2893 VSS.n1517 VSS.n313 3.32459
R2894 VSS.n1513 VSS.n312 3.32459
R2895 VSS.n1508 VSS.n311 3.32459
R2896 VSS.n1504 VSS.n310 3.32459
R2897 VSS.n1500 VSS.n309 3.32459
R2898 VSS.n1496 VSS.n308 3.32459
R2899 VSS.n1494 VSS.n319 3.32459
R2900 VSS.n614 VSS.n613 3.32459
R2901 VSS.n609 VSS.n607 3.32459
R2902 VSS.n622 VSS.n621 3.32459
R2903 VSS.n606 VSS.n604 3.32459
R2904 VSS.n629 VSS.n628 3.32459
R2905 VSS.n660 VSS.n655 3.32459
R2906 VSS.n663 VSS.n656 3.32459
R2907 VSS.n699 VSS.n698 3.32459
R2908 VSS.n679 VSS.n463 3.32459
R2909 VSS.n675 VSS.n464 3.32459
R2910 VSS.n1205 VSS.n465 3.32459
R2911 VSS.n467 VSS.n466 3.32459
R2912 VSS.n1210 VSS.n461 3.32459
R2913 VSS.n1212 VSS.n459 3.32459
R2914 VSS.n1233 VSS.n448 3.32459
R2915 VSS.n1238 VSS.n1237 3.32459
R2916 VSS.n1399 VSS.n386 3.32459
R2917 VSS.n1243 VSS.n1239 3.32459
R2918 VSS.n1246 VSS.n1240 3.32459
R2919 VSS.n1394 VSS.n1393 3.32459
R2920 VSS.n1264 VSS.n1263 3.32459
R2921 VSS.n1265 VSS.n1259 3.32459
R2922 VSS.n1272 VSS.n1271 3.32459
R2923 VSS.n1314 VSS.n1313 3.32459
R2924 VSS.n1309 VSS.n1275 3.32459
R2925 VSS.n1307 VSS.n1306 3.32459
R2926 VSS.n1287 VSS.n359 3.32459
R2927 VSS.n1283 VSS.n360 3.32459
R2928 VSS.n362 VSS.n361 3.32459
R2929 VSS.n369 VSS.n364 3.32459
R2930 VSS.n372 VSS.n365 3.32459
R2931 VSS.n1438 VSS.n1437 3.32459
R2932 VSS.n1418 VSS.n161 3.32459
R2933 VSS.n1414 VSS.n162 3.32459
R2934 VSS.n1951 VSS.n163 3.32459
R2935 VSS.n165 VSS.n164 3.32459
R2936 VSS.n1956 VSS.n159 3.32459
R2937 VSS.n1958 VSS.n157 3.32459
R2938 VSS.n1979 VSS.n146 3.32459
R2939 VSS.n1984 VSS.n1983 3.32459
R2940 VSS.n2013 VSS.n2011 3.32459
R2941 VSS.n1986 VSS.n1985 3.32459
R2942 VSS.n2009 VSS.n2008 3.32459
R2943 VSS.n2004 VSS.n1991 3.32459
R2944 VSS.n2289 VSS.n65 3.32459
R2945 VSS.n64 VSS.n58 3.32459
R2946 VSS.n2236 VSS.n63 3.32459
R2947 VSS.n2239 VSS.n61 3.32459
R2948 VSS.n2248 VSS.n50 3.32459
R2949 VSS.n2300 VSS.n2299 3.32459
R2950 VSS.n2300 VSS.n51 3.32459
R2951 VSS.n2247 VSS.n50 3.32459
R2952 VSS.n2237 VSS.n61 3.32459
R2953 VSS.n63 VSS.n62 3.32459
R2954 VSS.n2288 VSS.n64 3.32459
R2955 VSS.n67 VSS.n65 3.32459
R2956 VSS.n1991 VSS.n1988 3.32459
R2957 VSS.n2009 VSS.n1987 3.32459
R2958 VSS.n1985 VSS.n142 3.32459
R2959 VSS.n2011 VSS.n144 3.32459
R2960 VSS.n1984 VSS.n147 3.32459
R2961 VSS.n1977 VSS.n146 3.32459
R2962 VSS.n1959 VSS.n1958 3.32459
R2963 VSS.n1956 VSS.n1955 3.32459
R2964 VSS.n168 VSS.n164 3.32459
R2965 VSS.n1413 VSS.n163 3.32459
R2966 VSS.n1417 VSS.n162 3.32459
R2967 VSS.n1421 VSS.n161 3.32459
R2968 VSS.n1438 VSS.n366 3.32459
R2969 VSS.n370 VSS.n365 3.32459
R2970 VSS.n364 VSS.n363 3.32459
R2971 VSS.n1282 VSS.n362 3.32459
R2972 VSS.n1286 VSS.n360 3.32459
R2973 VSS.n1290 VSS.n359 3.32459
R2974 VSS.n1308 VSS.n1307 3.32459
R2975 VSS.n1275 VSS.n1273 3.32459
R2976 VSS.n1315 VSS.n1314 3.32459
R2977 VSS.n1271 VSS.n1270 3.32459
R2978 VSS.n1266 VSS.n1265 3.32459
R2979 VSS.n1263 VSS.n1262 3.32459
R2980 VSS.n1394 VSS.n1241 3.32459
R2981 VSS.n1244 VSS.n1240 3.32459
R2982 VSS.n1239 VSS.n385 3.32459
R2983 VSS.n450 VSS.n386 3.32459
R2984 VSS.n1238 VSS.n449 3.32459
R2985 VSS.n1231 VSS.n448 3.32459
R2986 VSS.n1213 VSS.n1212 3.32459
R2987 VSS.n1210 VSS.n1209 3.32459
R2988 VSS.n470 VSS.n466 3.32459
R2989 VSS.n674 VSS.n465 3.32459
R2990 VSS.n678 VSS.n464 3.32459
R2991 VSS.n682 VSS.n463 3.32459
R2992 VSS.n699 VSS.n657 3.32459
R2993 VSS.n661 VSS.n656 3.32459
R2994 VSS.n655 VSS.n653 3.32459
R2995 VSS.n2148 VSS.n2147 3.32459
R2996 VSS.n2149 VSS.n2144 3.32459
R2997 VSS.n2156 VSS.n2155 3.32459
R2998 VSS.n2157 VSS.n2141 3.32459
R2999 VSS.n2158 VSS.n2157 3.32459
R3000 VSS.n2155 VSS.n2154 3.32459
R3001 VSS.n2150 VSS.n2149 3.32459
R3002 VSS.n2147 VSS.n2146 3.32459
R3003 VSS.n2070 VSS.n10 2.53264
R3004 VSS.n2172 VSS.n2169 1.95679
R3005 VSS.n2298 VSS.n2297 1.4552
R3006 VSS VSS.n491 1.33138
R3007 VSS.n110 VSS.n1 1.32688
R3008 VSS.n1740 VSS.n1731 1.316
R3009 VSS.n1726 VSS.n233 1.316
R3010 VSS.n1007 VSS.n995 1.316
R3011 VSS.n973 VSS.n956 1.316
R3012 VSS.n906 VSS.n889 1.316
R3013 VSS.n838 VSS.n491 1.316
R3014 VSS.n810 VSS.n490 0.939203
R3015 VSS.n773 VSS.n490 0.939203
R3016 VSS.n803 VSS.n490 0.939203
R3017 VSS.n797 VSS.n490 0.939203
R3018 VSS.n795 VSS.n490 0.939203
R3019 VSS.n789 VSS.n490 0.939203
R3020 VSS.n787 VSS.n490 0.939203
R3021 VSS.n781 VSS.n490 0.939203
R3022 VSS.n814 VSS.n490 0.939203
R3023 VSS.n818 VSS.n490 0.939203
R3024 VSS.n2139 VSS.n97 0.939203
R3025 VSS.n2139 VSS.n95 0.939203
R3026 VSS.n2139 VSS.n94 0.939203
R3027 VSS.n2139 VSS.n93 0.939203
R3028 VSS.n2383 VSS.n3 0.939203
R3029 VSS.n2383 VSS.n4 0.939203
R3030 VSS.n114 VSS.n107 0.939203
R3031 VSS.n2101 VSS.n107 0.939203
R3032 VSS.n1738 VSS.n107 0.939203
R3033 VSS.n1744 VSS.n107 0.939203
R3034 VSS.n1736 VSS.n107 0.939203
R3035 VSS.n1751 VSS.n107 0.939203
R3036 VSS.n2056 VSS.n121 0.939203
R3037 VSS.n2056 VSS.n120 0.939203
R3038 VSS.n2056 VSS.n119 0.939203
R3039 VSS.n1765 VSS.n118 0.939203
R3040 VSS.n1772 VSS.n118 0.939203
R3041 VSS.n232 VSS.n118 0.939203
R3042 VSS.n1722 VSS.n118 0.939203
R3043 VSS.n1716 VSS.n118 0.939203
R3044 VSS.n1714 VSS.n222 0.939203
R3045 VSS.n1708 VSS.n1707 0.939203
R3046 VSS.n1699 VSS.n239 0.939203
R3047 VSS.n1700 VSS.n1699 0.939203
R3048 VSS.n1699 VSS.n254 0.939203
R3049 VSS.n1699 VSS.n246 0.939203
R3050 VSS.n1699 VSS.n245 0.939203
R3051 VSS.n1699 VSS.n244 0.939203
R3052 VSS.n1699 VSS.n243 0.939203
R3053 VSS.n1699 VSS.n242 0.939203
R3054 VSS.n1024 VSS.n1023 0.939203
R3055 VSS.n1001 VSS.n968 0.939203
R3056 VSS.n1031 VSS.n968 0.939203
R3057 VSS.n998 VSS.n968 0.939203
R3058 VSS.n1038 VSS.n968 0.939203
R3059 VSS.n1044 VSS.n968 0.939203
R3060 VSS.n971 VSS.n968 0.939203
R3061 VSS.n1051 VSS.n968 0.939203
R3062 VSS.n968 VSS.n967 0.939203
R3063 VSS.n1059 VSS.n1058 0.939203
R3064 VSS.n962 VSS.n901 0.939203
R3065 VSS.n1066 VSS.n901 0.939203
R3066 VSS.n959 VSS.n901 0.939203
R3067 VSS.n1073 VSS.n901 0.939203
R3068 VSS.n1079 VSS.n901 0.939203
R3069 VSS.n904 VSS.n901 0.939203
R3070 VSS.n1086 VSS.n901 0.939203
R3071 VSS.n901 VSS.n900 0.939203
R3072 VSS.n1094 VSS.n1093 0.939203
R3073 VSS.n895 VSS.n833 0.939203
R3074 VSS.n1101 VSS.n833 0.939203
R3075 VSS.n892 VSS.n833 0.939203
R3076 VSS.n1108 VSS.n833 0.939203
R3077 VSS.n1114 VSS.n833 0.939203
R3078 VSS.n836 VSS.n833 0.939203
R3079 VSS.n1121 VSS.n833 0.939203
R3080 VSS.n833 VSS.n832 0.939203
R3081 VSS.n1129 VSS.n1128 0.939203
R3082 VSS.n555 VSS.n545 0.939203
R3083 VSS.n549 VSS.n545 0.939203
R3084 VSS.n562 VSS.n545 0.939203
R3085 VSS.n565 VSS.n545 0.939203
R3086 VSS.n27 VSS.n24 0.939203
R3087 VSS.n2206 VSS.n27 0.939203
R3088 VSS.n2213 VSS.n27 0.939203
R3089 VSS.n2029 VSS.n2028 0.939203
R3090 VSS.n2028 VSS.n129 0.939203
R3091 VSS.n1864 VSS.n207 0.939203
R3092 VSS.n1867 VSS.n207 0.939203
R3093 VSS.n1873 VSS.n207 0.939203
R3094 VSS.n210 VSS.n207 0.939203
R3095 VSS.n1880 VSS.n207 0.939203
R3096 VSS.n223 VSS.n206 0.939203
R3097 VSS.n1888 VSS.n1887 0.939203
R3098 VSS.n201 VSS.n195 0.939203
R3099 VSS.n1895 VSS.n195 0.939203
R3100 VSS.n198 VSS.n195 0.939203
R3101 VSS.n1902 VSS.n195 0.939203
R3102 VSS.n1600 VSS.n195 0.939203
R3103 VSS.n1606 VSS.n195 0.939203
R3104 VSS.n1599 VSS.n195 0.939203
R3105 VSS.n1613 VSS.n195 0.939203
R3106 VSS.n1616 VSS.n1595 0.939203
R3107 VSS.n1622 VSS.n279 0.939203
R3108 VSS.n1592 VSS.n279 0.939203
R3109 VSS.n1629 VSS.n279 0.939203
R3110 VSS.n1632 VSS.n279 0.939203
R3111 VSS.n1585 VSS.n279 0.939203
R3112 VSS.n283 VSS.n279 0.939203
R3113 VSS.n1578 VSS.n279 0.939203
R3114 VSS.n1572 VSS.n279 0.939203
R3115 VSS.n1570 VSS.n1569 0.939203
R3116 VSS.n1562 VSS.n1561 0.939203
R3117 VSS.n1561 VSS.n1560 0.939203
R3118 VSS.n1561 VSS.n297 0.939203
R3119 VSS.n1561 VSS.n296 0.939203
R3120 VSS.n1561 VSS.n295 0.939203
R3121 VSS.n1561 VSS.n294 0.939203
R3122 VSS.n1561 VSS.n293 0.939203
R3123 VSS.n1561 VSS.n292 0.939203
R3124 VSS.n1532 VSS.n1531 0.939203
R3125 VSS.n1524 VSS.n1523 0.939203
R3126 VSS.n1523 VSS.n1522 0.939203
R3127 VSS.n1523 VSS.n313 0.939203
R3128 VSS.n1523 VSS.n312 0.939203
R3129 VSS.n1523 VSS.n311 0.939203
R3130 VSS.n1523 VSS.n310 0.939203
R3131 VSS.n1523 VSS.n309 0.939203
R3132 VSS.n1523 VSS.n308 0.939203
R3133 VSS.n1494 VSS.n1493 0.939203
R3134 VSS.n613 VSS.n521 0.939203
R3135 VSS.n609 VSS.n519 0.939203
R3136 VSS.n621 VSS.n519 0.939203
R3137 VSS.n606 VSS.n519 0.939203
R3138 VSS.n628 VSS.n519 0.939203
R3139 VSS.n2301 VSS.n2300 0.939203
R3140 VSS.n2301 VSS.n50 0.939203
R3141 VSS.n2294 VSS.n61 0.939203
R3142 VSS.n2294 VSS.n63 0.939203
R3143 VSS.n2294 VSS.n64 0.939203
R3144 VSS.n2294 VSS.n65 0.939203
R3145 VSS.n2010 VSS.n2009 0.939203
R3146 VSS.n2010 VSS.n1985 0.939203
R3147 VSS.n2011 VSS.n2010 0.939203
R3148 VSS.n2010 VSS.n1984 0.939203
R3149 VSS.n2010 VSS.n146 0.939203
R3150 VSS.n1958 VSS.n1957 0.939203
R3151 VSS.n1957 VSS.n1956 0.939203
R3152 VSS.n1957 VSS.n164 0.939203
R3153 VSS.n1957 VSS.n163 0.939203
R3154 VSS.n1957 VSS.n162 0.939203
R3155 VSS.n1957 VSS.n161 0.939203
R3156 VSS.n1439 VSS.n1438 0.939203
R3157 VSS.n1439 VSS.n365 0.939203
R3158 VSS.n1439 VSS.n364 0.939203
R3159 VSS.n1439 VSS.n362 0.939203
R3160 VSS.n1439 VSS.n360 0.939203
R3161 VSS.n1439 VSS.n359 0.939203
R3162 VSS.n1307 VSS.n1257 0.939203
R3163 VSS.n1275 VSS.n1257 0.939203
R3164 VSS.n1314 VSS.n1257 0.939203
R3165 VSS.n1271 VSS.n1257 0.939203
R3166 VSS.n1265 VSS.n1257 0.939203
R3167 VSS.n1263 VSS.n1257 0.939203
R3168 VSS.n1395 VSS.n1394 0.939203
R3169 VSS.n1395 VSS.n1240 0.939203
R3170 VSS.n1395 VSS.n1239 0.939203
R3171 VSS.n1395 VSS.n386 0.939203
R3172 VSS.n1395 VSS.n1238 0.939203
R3173 VSS.n1395 VSS.n448 0.939203
R3174 VSS.n1212 VSS.n1211 0.939203
R3175 VSS.n1211 VSS.n1210 0.939203
R3176 VSS.n1211 VSS.n466 0.939203
R3177 VSS.n1211 VSS.n465 0.939203
R3178 VSS.n1211 VSS.n464 0.939203
R3179 VSS.n1211 VSS.n463 0.939203
R3180 VSS.n700 VSS.n699 0.939203
R3181 VSS.n700 VSS.n656 0.939203
R3182 VSS.n700 VSS.n655 0.939203
R3183 VSS.n2157 VSS.n2139 0.939203
R3184 VSS.n2155 VSS.n2139 0.939203
R3185 VSS.n2149 VSS.n2139 0.939203
R3186 VSS.n2147 VSS.n2139 0.939203
R3187 VSS.n1997 VSS.n1996 0.931463
R3188 VSS.n2167 VSS.t3 0.8195
R3189 VSS.n2167 VSS.t15 0.8195
R3190 VSS.n2168 VSS.t7 0.8195
R3191 VSS.n2168 VSS.t10 0.8195
R3192 VSS.n154 VSS.n143 0.702875
R3193 VSS.n1406 VSS.n169 0.702875
R3194 VSS.n1405 VSS.n1404 0.702875
R3195 VSS.n1403 VSS.n1402 0.702875
R3196 VSS.n1401 VSS.n381 0.702875
R3197 VSS.n667 VSS.n471 0.702875
R3198 VSS.n1222 VSS.n456 0.698622
R3199 VSS.n377 VSS.n376 0.698622
R3200 VSS.n1968 VSS.n153 0.698622
R3201 VSS.n1407 VSS.n375 0.698622
R3202 VSS.n380 VSS.n379 0.698622
R3203 VSS.n668 VSS.n666 0.698622
R3204 VSS.n143 VSS.n53 0.692375
R3205 VSS.n667 VSS 0.629
R3206 VSS.n2297 VSS.n53 0.624125
R3207 VSS.n169 VSS.n154 0.613625
R3208 VSS.n1406 VSS.n1405 0.613625
R3209 VSS.n1404 VSS.n1403 0.613625
R3210 VSS.n1402 VSS.n1401 0.613625
R3211 VSS.n471 VSS.n381 0.613625
R3212 VSS VSS.n2385 0.397167
R3213 VSS.n2385 VSS.n1 0.367833
R3214 VSS.n662 VSS.n659 0.237342
R3215 VSS.n664 VSS.n662 0.237342
R3216 VSS.n665 VSS.n664 0.237342
R3217 VSS.n697 VSS.n665 0.237342
R3218 VSS.n697 VSS.n696 0.237342
R3219 VSS.n696 VSS.n695 0.237342
R3220 VSS.n689 VSS.n688 0.237342
R3221 VSS.n688 VSS.n687 0.237342
R3222 VSS.n687 VSS.n673 0.237342
R3223 VSS.n681 VSS.n673 0.237342
R3224 VSS.n681 VSS.n680 0.237342
R3225 VSS.n680 VSS.n677 0.237342
R3226 VSS.n677 VSS.n676 0.237342
R3227 VSS.n676 VSS.n468 0.237342
R3228 VSS.n1208 VSS.n1207 0.237342
R3229 VSS.n1208 VSS.n460 0.237342
R3230 VSS.n1214 VSS.n460 0.237342
R3231 VSS.n1215 VSS.n1214 0.237342
R3232 VSS.n1216 VSS.n1215 0.237342
R3233 VSS.n1216 VSS.n455 0.237342
R3234 VSS.n1225 VSS.n1223 0.237342
R3235 VSS.n1225 VSS.n1224 0.237342
R3236 VSS.n1224 VSS.n451 0.237342
R3237 VSS.n1232 VSS.n451 0.237342
R3238 VSS.n1234 VSS.n1232 0.237342
R3239 VSS.n1235 VSS.n1234 0.237342
R3240 VSS.n1236 VSS.n1235 0.237342
R3241 VSS.n1236 VSS.n382 0.237342
R3242 VSS.n1245 VSS.n383 0.237342
R3243 VSS.n1247 VSS.n1245 0.237342
R3244 VSS.n1248 VSS.n1247 0.237342
R3245 VSS.n1392 VSS.n1248 0.237342
R3246 VSS.n1392 VSS.n1391 0.237342
R3247 VSS.n1391 VSS.n1390 0.237342
R3248 VSS.n1384 VSS.n1383 0.237342
R3249 VSS.n1383 VSS.n1382 0.237342
R3250 VSS.n1382 VSS.n1253 0.237342
R3251 VSS.n1261 VSS.n1253 0.237342
R3252 VSS.n1261 VSS.n1260 0.237342
R3253 VSS.n1267 VSS.n1260 0.237342
R3254 VSS.n1268 VSS.n1267 0.237342
R3255 VSS.n1269 VSS.n1268 0.237342
R3256 VSS.n1312 VSS.n1311 0.237342
R3257 VSS.n1311 VSS.n1310 0.237342
R3258 VSS.n1310 VSS.n1274 0.237342
R3259 VSS.n1305 VSS.n1274 0.237342
R3260 VSS.n1305 VSS.n1304 0.237342
R3261 VSS.n1304 VSS.n1303 0.237342
R3262 VSS.n1297 VSS.n1296 0.237342
R3263 VSS.n1296 VSS.n1295 0.237342
R3264 VSS.n1295 VSS.n1280 0.237342
R3265 VSS.n1289 VSS.n1280 0.237342
R3266 VSS.n1289 VSS.n1288 0.237342
R3267 VSS.n1288 VSS.n1285 0.237342
R3268 VSS.n1285 VSS.n1284 0.237342
R3269 VSS.n1284 VSS.n1281 0.237342
R3270 VSS.n371 VSS.n368 0.237342
R3271 VSS.n373 VSS.n371 0.237342
R3272 VSS.n374 VSS.n373 0.237342
R3273 VSS.n1436 VSS.n374 0.237342
R3274 VSS.n1436 VSS.n1435 0.237342
R3275 VSS.n1435 VSS.n1434 0.237342
R3276 VSS.n1428 VSS.n1427 0.237342
R3277 VSS.n1427 VSS.n1426 0.237342
R3278 VSS.n1426 VSS.n1412 0.237342
R3279 VSS.n1420 VSS.n1412 0.237342
R3280 VSS.n1420 VSS.n1419 0.237342
R3281 VSS.n1419 VSS.n1416 0.237342
R3282 VSS.n1416 VSS.n1415 0.237342
R3283 VSS.n1415 VSS.n166 0.237342
R3284 VSS.n1954 VSS.n1953 0.237342
R3285 VSS.n1954 VSS.n158 0.237342
R3286 VSS.n1960 VSS.n158 0.237342
R3287 VSS.n1961 VSS.n1960 0.237342
R3288 VSS.n1962 VSS.n1961 0.237342
R3289 VSS.n1962 VSS.n152 0.237342
R3290 VSS.n1971 VSS.n1969 0.237342
R3291 VSS.n1971 VSS.n1970 0.237342
R3292 VSS.n1970 VSS.n148 0.237342
R3293 VSS.n1978 VSS.n148 0.237342
R3294 VSS.n1980 VSS.n1978 0.237342
R3295 VSS.n1981 VSS.n1980 0.237342
R3296 VSS.n1982 VSS.n1981 0.237342
R3297 VSS.n1982 VSS.n140 0.237342
R3298 VSS.n1989 VSS.n141 0.237342
R3299 VSS.n2007 VSS.n1989 0.237342
R3300 VSS.n2007 VSS.n2006 0.237342
R3301 VSS.n2006 VSS.n2005 0.237342
R3302 VSS.n2005 VSS.n1990 0.237342
R3303 VSS.n1995 VSS.n1990 0.237342
R3304 VSS.n1998 VSS.n1995 0.237342
R3305 VSS.n2285 VSS.n68 0.237342
R3306 VSS.n2286 VSS.n2285 0.237342
R3307 VSS.n2292 VSS.n2286 0.237342
R3308 VSS.n2292 VSS.n2291 0.237342
R3309 VSS.n2291 VSS.n2290 0.237342
R3310 VSS.n2290 VSS.n2287 0.237342
R3311 VSS.n2287 VSS.n54 0.237342
R3312 VSS.n2235 VSS.n55 0.237342
R3313 VSS.n2238 VSS.n2235 0.237342
R3314 VSS.n2240 VSS.n2238 0.237342
R3315 VSS.n2241 VSS.n2240 0.237342
R3316 VSS.n2267 VSS.n2241 0.237342
R3317 VSS.n2267 VSS.n2266 0.237342
R3318 VSS.n2266 VSS.n2265 0.237342
R3319 VSS.n2265 VSS.n2242 0.237342
R3320 VSS.n2259 VSS.n2242 0.237342
R3321 VSS.n2259 VSS.n2258 0.237342
R3322 VSS.n2258 VSS.n2257 0.237342
R3323 VSS.n2257 VSS.n2246 0.237342
R3324 VSS.n2251 VSS.n2246 0.237342
R3325 VSS.n2251 VSS.n2250 0.237342
R3326 VSS.n2250 VSS.n2249 0.237342
R3327 VSS.n2249 VSS.n52 0.237342
R3328 VSS.n546 VSS.n544 0.237342
R3329 VSS.n560 VSS.n546 0.237342
R3330 VSS.n560 VSS.n559 0.237342
R3331 VSS.n559 VSS.n558 0.237342
R3332 VSS.n558 VSS.n548 0.237342
R3333 VSS.n553 VSS.n548 0.237342
R3334 VSS.n553 VSS.n552 0.237342
R3335 VSS.n552 VSS.n515 0.237342
R3336 VSS.n747 VSS.n515 0.237342
R3337 VSS.n748 VSS.n747 0.237342
R3338 VSS.n749 VSS.n748 0.237342
R3339 VSS.n749 VSS.n506 0.237342
R3340 VSS.n762 VSS.n506 0.237342
R3341 VSS.n763 VSS.n762 0.237342
R3342 VSS.n764 VSS.n763 0.237342
R3343 VSS.n764 VSS.n495 0.237342
R3344 VSS.n2145 VSS.n87 0.237342
R3345 VSS.n2151 VSS.n2145 0.237342
R3346 VSS.n2152 VSS.n2151 0.237342
R3347 VSS.n2153 VSS.n2152 0.237342
R3348 VSS.n2153 VSS.n2143 0.237342
R3349 VSS.n2159 VSS.n2143 0.237342
R3350 VSS.n2160 VSS.n2159 0.237342
R3351 VSS.n2182 VSS.n2160 0.237342
R3352 VSS.n2182 VSS.n2181 0.237342
R3353 VSS.n2181 VSS.n2180 0.237342
R3354 VSS.n2180 VSS.n2161 0.237342
R3355 VSS.n2174 VSS.n2161 0.237342
R3356 VSS.n2174 VSS.n2173 0.237342
R3357 VSS.n2315 VSS.n2314 0.237342
R3358 VSS.n2314 VSS.n43 0.237342
R3359 VSS.n2308 VSS.n43 0.237342
R3360 VSS.n2308 VSS.n2307 0.237342
R3361 VSS.n2307 VSS.n2306 0.237342
R3362 VSS.n2306 VSS.n47 0.237342
R3363 VSS.n2330 VSS.n35 0.237342
R3364 VSS.n2324 VSS.n35 0.237342
R3365 VSS.n2324 VSS.n2323 0.237342
R3366 VSS.n2323 VSS.n2322 0.237342
R3367 VSS.n2322 VSS.n39 0.237342
R3368 VSS.n2099 VSS.n111 0.237342
R3369 VSS.n2099 VSS.n2098 0.237342
R3370 VSS.n2098 VSS.n2097 0.237342
R3371 VSS.n2097 VSS.n113 0.237342
R3372 VSS.n2061 VSS.n113 0.237342
R3373 VSS.n2090 VSS.n2061 0.237342
R3374 VSS.n2090 VSS.n2089 0.237342
R3375 VSS.n2089 VSS.n2088 0.237342
R3376 VSS.n2088 VSS.n2062 0.237342
R3377 VSS.n2082 VSS.n2062 0.237342
R3378 VSS.n2082 VSS.n2081 0.237342
R3379 VSS.n2081 VSS.n2080 0.237342
R3380 VSS.n2080 VSS.n2066 0.237342
R3381 VSS.n2074 VSS.n2066 0.237342
R3382 VSS.n2074 VSS.n2073 0.237342
R3383 VSS.n2073 VSS.n2072 0.237342
R3384 VSS.n1150 VSS.n496 0.237342
R3385 VSS.n1150 VSS.n1149 0.237342
R3386 VSS.n1149 VSS.n1148 0.237342
R3387 VSS.n1148 VSS.n826 0.237342
R3388 VSS.n1133 VSS.n826 0.237342
R3389 VSS.n1133 VSS.n1132 0.237342
R3390 VSS.n1132 VSS.n1131 0.237342
R3391 VSS.n1131 VSS.n828 0.237342
R3392 VSS.n1126 VSS.n828 0.237342
R3393 VSS.n1126 VSS.n1125 0.237342
R3394 VSS.n1125 VSS.n1124 0.237342
R3395 VSS.n1124 VSS.n831 0.237342
R3396 VSS.n1119 VSS.n831 0.237342
R3397 VSS.n1119 VSS.n1118 0.237342
R3398 VSS.n1118 VSS.n1117 0.237342
R3399 VSS.n1117 VSS.n835 0.237342
R3400 VSS.n2106 VSS.n105 0.237342
R3401 VSS.n2112 VSS.n105 0.237342
R3402 VSS.n2113 VSS.n2112 0.237342
R3403 VSS.n2114 VSS.n2113 0.237342
R3404 VSS.n2114 VSS.n101 0.237342
R3405 VSS.n2120 VSS.n101 0.237342
R3406 VSS.n2121 VSS.n2120 0.237342
R3407 VSS.n2135 VSS.n2121 0.237342
R3408 VSS.n2135 VSS.n2134 0.237342
R3409 VSS.n2134 VSS.n2133 0.237342
R3410 VSS.n2133 VSS.n2130 0.237342
R3411 VSS.n2130 VSS.n2129 0.237342
R3412 VSS.n2129 VSS.n2126 0.237342
R3413 VSS.n2126 VSS.n2125 0.237342
R3414 VSS.n2125 VSS.n2122 0.237342
R3415 VSS.n2122 VSS.n88 0.237342
R3416 VSS.n1770 VSS.n1769 0.237342
R3417 VSS.n1769 VSS.n1768 0.237342
R3418 VSS.n1768 VSS.n1764 0.237342
R3419 VSS.n1764 VSS.n1763 0.237342
R3420 VSS.n1763 VSS.n1760 0.237342
R3421 VSS.n1760 VSS.n1759 0.237342
R3422 VSS.n1759 VSS.n1756 0.237342
R3423 VSS.n1756 VSS.n1755 0.237342
R3424 VSS.n1755 VSS.n1732 0.237342
R3425 VSS.n1733 VSS.n1732 0.237342
R3426 VSS.n1749 VSS.n1733 0.237342
R3427 VSS.n1749 VSS.n1748 0.237342
R3428 VSS.n1748 VSS.n1747 0.237342
R3429 VSS.n1747 VSS.n1735 0.237342
R3430 VSS.n1742 VSS.n1735 0.237342
R3431 VSS.n1742 VSS.n1741 0.237342
R3432 VSS.n1778 VSS.n1777 0.237342
R3433 VSS.n1779 VSS.n1778 0.237342
R3434 VSS.n1779 VSS.n227 0.237342
R3435 VSS.n1785 VSS.n227 0.237342
R3436 VSS.n1786 VSS.n1785 0.237342
R3437 VSS.n1787 VSS.n1786 0.237342
R3438 VSS.n1787 VSS.n220 0.237342
R3439 VSS.n1794 VSS.n220 0.237342
R3440 VSS.n1795 VSS.n1794 0.237342
R3441 VSS.n1796 VSS.n1795 0.237342
R3442 VSS.n1796 VSS.n216 0.237342
R3443 VSS.n1802 VSS.n216 0.237342
R3444 VSS.n1803 VSS.n1802 0.237342
R3445 VSS.n1804 VSS.n1803 0.237342
R3446 VSS.n1804 VSS.n212 0.237342
R3447 VSS.n1810 VSS.n212 0.237342
R3448 VSS.n250 VSS.n249 0.237342
R3449 VSS.n252 VSS.n250 0.237342
R3450 VSS.n252 VSS.n251 0.237342
R3451 VSS.n251 VSS.n240 0.237342
R3452 VSS.n1703 VSS.n240 0.237342
R3453 VSS.n1704 VSS.n1703 0.237342
R3454 VSS.n1704 VSS.n238 0.237342
R3455 VSS.n1710 VSS.n238 0.237342
R3456 VSS.n1711 VSS.n1710 0.237342
R3457 VSS.n1712 VSS.n1711 0.237342
R3458 VSS.n1712 VSS.n236 0.237342
R3459 VSS.n1718 VSS.n236 0.237342
R3460 VSS.n1719 VSS.n1718 0.237342
R3461 VSS.n1720 VSS.n1719 0.237342
R3462 VSS.n1720 VSS.n234 0.237342
R3463 VSS.n1725 VSS.n234 0.237342
R3464 VSS.n1696 VSS.n1695 0.237342
R3465 VSS.n1695 VSS.n1694 0.237342
R3466 VSS.n1694 VSS.n261 0.237342
R3467 VSS.n1688 VSS.n261 0.237342
R3468 VSS.n1688 VSS.n1687 0.237342
R3469 VSS.n1687 VSS.n1686 0.237342
R3470 VSS.n1686 VSS.n265 0.237342
R3471 VSS.n1679 VSS.n265 0.237342
R3472 VSS.n1679 VSS.n1678 0.237342
R3473 VSS.n1678 VSS.n1677 0.237342
R3474 VSS.n1677 VSS.n1658 0.237342
R3475 VSS.n1671 VSS.n1658 0.237342
R3476 VSS.n1671 VSS.n1670 0.237342
R3477 VSS.n1670 VSS.n1669 0.237342
R3478 VSS.n1669 VSS.n1663 0.237342
R3479 VSS.n1663 VSS.n1662 0.237342
R3480 VSS.n1036 VSS.n1035 0.237342
R3481 VSS.n1035 VSS.n1034 0.237342
R3482 VSS.n1034 VSS.n997 0.237342
R3483 VSS.n1029 VSS.n997 0.237342
R3484 VSS.n1029 VSS.n1028 0.237342
R3485 VSS.n1028 VSS.n1027 0.237342
R3486 VSS.n1027 VSS.n1000 0.237342
R3487 VSS.n1004 VSS.n1000 0.237342
R3488 VSS.n1021 VSS.n1004 0.237342
R3489 VSS.n1021 VSS.n1020 0.237342
R3490 VSS.n1020 VSS.n1019 0.237342
R3491 VSS.n1019 VSS.n1016 0.237342
R3492 VSS.n1016 VSS.n1015 0.237342
R3493 VSS.n1015 VSS.n1012 0.237342
R3494 VSS.n1012 VSS.n1011 0.237342
R3495 VSS.n1011 VSS.n1008 0.237342
R3496 VSS.n994 VSS.n974 0.237342
R3497 VSS.n988 VSS.n974 0.237342
R3498 VSS.n988 VSS.n987 0.237342
R3499 VSS.n987 VSS.n986 0.237342
R3500 VSS.n986 VSS.n978 0.237342
R3501 VSS.n980 VSS.n978 0.237342
R3502 VSS.n980 VSS.n272 0.237342
R3503 VSS.n1652 VSS.n272 0.237342
R3504 VSS.n1652 VSS.n1651 0.237342
R3505 VSS.n1651 VSS.n1650 0.237342
R3506 VSS.n1650 VSS.n273 0.237342
R3507 VSS.n1644 VSS.n273 0.237342
R3508 VSS.n1644 VSS.n1643 0.237342
R3509 VSS.n1643 VSS.n1642 0.237342
R3510 VSS.n1642 VSS.n277 0.237342
R3511 VSS.n1636 VSS.n277 0.237342
R3512 VSS.n1071 VSS.n1070 0.237342
R3513 VSS.n1070 VSS.n1069 0.237342
R3514 VSS.n1069 VSS.n958 0.237342
R3515 VSS.n1064 VSS.n958 0.237342
R3516 VSS.n1064 VSS.n1063 0.237342
R3517 VSS.n1063 VSS.n1062 0.237342
R3518 VSS.n1062 VSS.n961 0.237342
R3519 VSS.n965 VSS.n961 0.237342
R3520 VSS.n1056 VSS.n965 0.237342
R3521 VSS.n1056 VSS.n1055 0.237342
R3522 VSS.n1055 VSS.n1054 0.237342
R3523 VSS.n1054 VSS.n966 0.237342
R3524 VSS.n1049 VSS.n966 0.237342
R3525 VSS.n1049 VSS.n1048 0.237342
R3526 VSS.n1048 VSS.n1047 0.237342
R3527 VSS.n1047 VSS.n970 0.237342
R3528 VSS.n955 VSS.n907 0.237342
R3529 VSS.n949 VSS.n907 0.237342
R3530 VSS.n949 VSS.n948 0.237342
R3531 VSS.n948 VSS.n947 0.237342
R3532 VSS.n947 VSS.n911 0.237342
R3533 VSS.n941 VSS.n911 0.237342
R3534 VSS.n941 VSS.n940 0.237342
R3535 VSS.n940 VSS.n939 0.237342
R3536 VSS.n939 VSS.n915 0.237342
R3537 VSS.n933 VSS.n915 0.237342
R3538 VSS.n933 VSS.n932 0.237342
R3539 VSS.n932 VSS.n931 0.237342
R3540 VSS.n931 VSS.n919 0.237342
R3541 VSS.n925 VSS.n919 0.237342
R3542 VSS.n925 VSS.n924 0.237342
R3543 VSS.n924 VSS.n923 0.237342
R3544 VSS.n1106 VSS.n1105 0.237342
R3545 VSS.n1105 VSS.n1104 0.237342
R3546 VSS.n1104 VSS.n891 0.237342
R3547 VSS.n1099 VSS.n891 0.237342
R3548 VSS.n1099 VSS.n1098 0.237342
R3549 VSS.n1098 VSS.n1097 0.237342
R3550 VSS.n1097 VSS.n894 0.237342
R3551 VSS.n898 VSS.n894 0.237342
R3552 VSS.n1091 VSS.n898 0.237342
R3553 VSS.n1091 VSS.n1090 0.237342
R3554 VSS.n1090 VSS.n1089 0.237342
R3555 VSS.n1089 VSS.n899 0.237342
R3556 VSS.n1084 VSS.n899 0.237342
R3557 VSS.n1084 VSS.n1083 0.237342
R3558 VSS.n1083 VSS.n1082 0.237342
R3559 VSS.n1082 VSS.n903 0.237342
R3560 VSS.n888 VSS.n839 0.237342
R3561 VSS.n882 VSS.n839 0.237342
R3562 VSS.n882 VSS.n881 0.237342
R3563 VSS.n881 VSS.n880 0.237342
R3564 VSS.n880 VSS.n843 0.237342
R3565 VSS.n874 VSS.n843 0.237342
R3566 VSS.n874 VSS.n873 0.237342
R3567 VSS.n873 VSS.n872 0.237342
R3568 VSS.n872 VSS.n847 0.237342
R3569 VSS.n866 VSS.n847 0.237342
R3570 VSS.n866 VSS.n865 0.237342
R3571 VSS.n865 VSS.n864 0.237342
R3572 VSS.n864 VSS.n852 0.237342
R3573 VSS.n858 VSS.n852 0.237342
R3574 VSS.n858 VSS.n857 0.237342
R3575 VSS.n857 VSS.n856 0.237342
R3576 VSS.n783 VSS.n497 0.237342
R3577 VSS.n784 VSS.n783 0.237342
R3578 VSS.n785 VSS.n784 0.237342
R3579 VSS.n785 VSS.n778 0.237342
R3580 VSS.n791 VSS.n778 0.237342
R3581 VSS.n792 VSS.n791 0.237342
R3582 VSS.n793 VSS.n792 0.237342
R3583 VSS.n793 VSS.n776 0.237342
R3584 VSS.n799 VSS.n776 0.237342
R3585 VSS.n800 VSS.n799 0.237342
R3586 VSS.n801 VSS.n800 0.237342
R3587 VSS.n801 VSS.n774 0.237342
R3588 VSS.n806 VSS.n774 0.237342
R3589 VSS.n807 VSS.n806 0.237342
R3590 VSS.n807 VSS.n772 0.237342
R3591 VSS.n812 VSS.n772 0.237342
R3592 VSS.n1855 VSS.n1811 0.237342
R3593 VSS.n1849 VSS.n1811 0.237342
R3594 VSS.n1849 VSS.n1848 0.237342
R3595 VSS.n1848 VSS.n1847 0.237342
R3596 VSS.n1847 VSS.n1815 0.237342
R3597 VSS.n1841 VSS.n1815 0.237342
R3598 VSS.n1841 VSS.n1840 0.237342
R3599 VSS.n1840 VSS.n1839 0.237342
R3600 VSS.n1839 VSS.n1819 0.237342
R3601 VSS.n1833 VSS.n1819 0.237342
R3602 VSS.n1833 VSS.n1832 0.237342
R3603 VSS.n1832 VSS.n1831 0.237342
R3604 VSS.n1831 VSS.n1823 0.237342
R3605 VSS.n1825 VSS.n1823 0.237342
R3606 VSS.n1825 VSS.n135 0.237342
R3607 VSS.n2024 VSS.n135 0.237342
R3608 VSS.n2024 VSS.n2023 0.237342
R3609 VSS.n2023 VSS.n2022 0.237342
R3610 VSS.n2022 VSS.n136 0.237342
R3611 VSS.n2016 VSS.n136 0.237342
R3612 VSS.n2016 VSS.n2015 0.237342
R3613 VSS.n1908 VSS.n1907 0.237342
R3614 VSS.n1909 VSS.n1908 0.237342
R3615 VSS.n1909 VSS.n186 0.237342
R3616 VSS.n1916 VSS.n186 0.237342
R3617 VSS.n1917 VSS.n1916 0.237342
R3618 VSS.n1918 VSS.n1917 0.237342
R3619 VSS.n1918 VSS.n182 0.237342
R3620 VSS.n1924 VSS.n182 0.237342
R3621 VSS.n1925 VSS.n1924 0.237342
R3622 VSS.n1926 VSS.n1925 0.237342
R3623 VSS.n1926 VSS.n178 0.237342
R3624 VSS.n1932 VSS.n178 0.237342
R3625 VSS.n1933 VSS.n1932 0.237342
R3626 VSS.n1934 VSS.n1933 0.237342
R3627 VSS.n1934 VSS.n174 0.237342
R3628 VSS.n1940 VSS.n174 0.237342
R3629 VSS.n1941 VSS.n1940 0.237342
R3630 VSS.n1943 VSS.n1941 0.237342
R3631 VSS.n1943 VSS.n1942 0.237342
R3632 VSS.n1942 VSS.n171 0.237342
R3633 VSS.n171 VSS.n167 0.237342
R3634 VSS.n338 VSS.n281 0.237342
R3635 VSS.n339 VSS.n338 0.237342
R3636 VSS.n1476 VSS.n339 0.237342
R3637 VSS.n1476 VSS.n1475 0.237342
R3638 VSS.n1475 VSS.n1474 0.237342
R3639 VSS.n1474 VSS.n340 0.237342
R3640 VSS.n1468 VSS.n340 0.237342
R3641 VSS.n1468 VSS.n1467 0.237342
R3642 VSS.n1467 VSS.n1466 0.237342
R3643 VSS.n1466 VSS.n344 0.237342
R3644 VSS.n1460 VSS.n344 0.237342
R3645 VSS.n1460 VSS.n1459 0.237342
R3646 VSS.n1459 VSS.n1458 0.237342
R3647 VSS.n1458 VSS.n348 0.237342
R3648 VSS.n1452 VSS.n348 0.237342
R3649 VSS.n1452 VSS.n1451 0.237342
R3650 VSS.n1451 VSS.n1450 0.237342
R3651 VSS.n1450 VSS.n352 0.237342
R3652 VSS.n1444 VSS.n352 0.237342
R3653 VSS.n1444 VSS.n1443 0.237342
R3654 VSS.n1443 VSS.n1442 0.237342
R3655 VSS.n1334 VSS.n1333 0.237342
R3656 VSS.n1334 VSS.n1332 0.237342
R3657 VSS.n1341 VSS.n1332 0.237342
R3658 VSS.n1342 VSS.n1341 0.237342
R3659 VSS.n1343 VSS.n1342 0.237342
R3660 VSS.n1343 VSS.n1329 0.237342
R3661 VSS.n1349 VSS.n1329 0.237342
R3662 VSS.n1350 VSS.n1349 0.237342
R3663 VSS.n1351 VSS.n1350 0.237342
R3664 VSS.n1351 VSS.n1325 0.237342
R3665 VSS.n1357 VSS.n1325 0.237342
R3666 VSS.n1358 VSS.n1357 0.237342
R3667 VSS.n1359 VSS.n1358 0.237342
R3668 VSS.n1359 VSS.n1321 0.237342
R3669 VSS.n1365 VSS.n1321 0.237342
R3670 VSS.n1366 VSS.n1365 0.237342
R3671 VSS.n1367 VSS.n1366 0.237342
R3672 VSS.n1367 VSS.n1317 0.237342
R3673 VSS.n1373 VSS.n1317 0.237342
R3674 VSS.n1374 VSS.n1373 0.237342
R3675 VSS.n1375 VSS.n1374 0.237342
R3676 VSS.n409 VSS.n404 0.237342
R3677 VSS.n410 VSS.n409 0.237342
R3678 VSS.n411 VSS.n410 0.237342
R3679 VSS.n411 VSS.n402 0.237342
R3680 VSS.n416 VSS.n402 0.237342
R3681 VSS.n417 VSS.n416 0.237342
R3682 VSS.n418 VSS.n417 0.237342
R3683 VSS.n418 VSS.n398 0.237342
R3684 VSS.n424 VSS.n398 0.237342
R3685 VSS.n425 VSS.n424 0.237342
R3686 VSS.n426 VSS.n425 0.237342
R3687 VSS.n426 VSS.n394 0.237342
R3688 VSS.n432 VSS.n394 0.237342
R3689 VSS.n433 VSS.n432 0.237342
R3690 VSS.n434 VSS.n433 0.237342
R3691 VSS.n434 VSS.n390 0.237342
R3692 VSS.n440 VSS.n390 0.237342
R3693 VSS.n441 VSS.n440 0.237342
R3694 VSS.n443 VSS.n441 0.237342
R3695 VSS.n443 VSS.n442 0.237342
R3696 VSS.n442 VSS.n384 0.237342
R3697 VSS.n820 VSS.n813 0.237342
R3698 VSS.n815 VSS.n813 0.237342
R3699 VSS.n815 VSS.n488 0.237342
R3700 VSS.n1170 VSS.n488 0.237342
R3701 VSS.n1171 VSS.n1170 0.237342
R3702 VSS.n1172 VSS.n1171 0.237342
R3703 VSS.n1172 VSS.n484 0.237342
R3704 VSS.n1178 VSS.n484 0.237342
R3705 VSS.n1179 VSS.n1178 0.237342
R3706 VSS.n1180 VSS.n1179 0.237342
R3707 VSS.n1180 VSS.n480 0.237342
R3708 VSS.n1186 VSS.n480 0.237342
R3709 VSS.n1187 VSS.n1186 0.237342
R3710 VSS.n1188 VSS.n1187 0.237342
R3711 VSS.n1188 VSS.n476 0.237342
R3712 VSS.n1194 VSS.n476 0.237342
R3713 VSS.n1195 VSS.n1194 0.237342
R3714 VSS.n1197 VSS.n1195 0.237342
R3715 VSS.n1197 VSS.n1196 0.237342
R3716 VSS.n1196 VSS.n473 0.237342
R3717 VSS.n473 VSS.n469 0.237342
R3718 VSS.n634 VSS.n526 0.237342
R3719 VSS.n635 VSS.n634 0.237342
R3720 VSS.n737 VSS.n635 0.237342
R3721 VSS.n737 VSS.n736 0.237342
R3722 VSS.n736 VSS.n735 0.237342
R3723 VSS.n735 VSS.n636 0.237342
R3724 VSS.n729 VSS.n636 0.237342
R3725 VSS.n729 VSS.n728 0.237342
R3726 VSS.n728 VSS.n727 0.237342
R3727 VSS.n727 VSS.n640 0.237342
R3728 VSS.n721 VSS.n640 0.237342
R3729 VSS.n721 VSS.n720 0.237342
R3730 VSS.n720 VSS.n719 0.237342
R3731 VSS.n719 VSS.n644 0.237342
R3732 VSS.n713 VSS.n644 0.237342
R3733 VSS.n713 VSS.n712 0.237342
R3734 VSS.n712 VSS.n711 0.237342
R3735 VSS.n711 VSS.n648 0.237342
R3736 VSS.n705 VSS.n648 0.237342
R3737 VSS.n705 VSS.n704 0.237342
R3738 VSS.n704 VSS.n703 0.237342
R3739 VSS.n2381 VSS.n2380 0.237342
R3740 VSS.n2380 VSS.n2379 0.237342
R3741 VSS.n2379 VSS.n2376 0.237342
R3742 VSS.n2376 VSS.n2375 0.237342
R3743 VSS.n2375 VSS.n8 0.237342
R3744 VSS.n13 VSS.n8 0.237342
R3745 VSS.n2368 VSS.n13 0.237342
R3746 VSS.n2366 VSS.n2365 0.237342
R3747 VSS.n2365 VSS.n14 0.237342
R3748 VSS.n2359 VSS.n14 0.237342
R3749 VSS.n2359 VSS.n2358 0.237342
R3750 VSS.n2358 VSS.n2357 0.237342
R3751 VSS.n2357 VSS.n18 0.237342
R3752 VSS.n2351 VSS.n18 0.237342
R3753 VSS.n2351 VSS.n2350 0.237342
R3754 VSS.n30 VSS.n22 0.237342
R3755 VSS.n2340 VSS.n30 0.237342
R3756 VSS.n2340 VSS.n2339 0.237342
R3757 VSS.n2339 VSS.n2338 0.237342
R3758 VSS.n2338 VSS.n31 0.237342
R3759 VSS.n2332 VSS.n31 0.237342
R3760 VSS.n626 VSS.n603 0.237342
R3761 VSS.n626 VSS.n625 0.237342
R3762 VSS.n625 VSS.n624 0.237342
R3763 VSS.n624 VSS.n605 0.237342
R3764 VSS.n619 VSS.n605 0.237342
R3765 VSS.n619 VSS.n618 0.237342
R3766 VSS.n618 VSS.n617 0.237342
R3767 VSS.n617 VSS.n608 0.237342
R3768 VSS.n610 VSS.n608 0.237342
R3769 VSS.n611 VSS.n610 0.237342
R3770 VSS.n611 VSS.n511 0.237342
R3771 VSS.n755 VSS.n511 0.237342
R3772 VSS.n756 VSS.n755 0.237342
R3773 VSS.n757 VSS.n756 0.237342
R3774 VSS.n757 VSS.n502 0.237342
R3775 VSS.n770 VSS.n502 0.237342
R3776 VSS.n771 VSS.n770 0.237342
R3777 VSS.n1158 VSS.n771 0.237342
R3778 VSS.n1156 VSS.n821 0.237342
R3779 VSS.n1141 VSS.n821 0.237342
R3780 VSS.n1142 VSS.n1141 0.237342
R3781 VSS.n1143 VSS.n1142 0.237342
R3782 VSS.n1143 VSS.n321 0.237342
R3783 VSS.n1488 VSS.n321 0.237342
R3784 VSS.n1489 VSS.n1488 0.237342
R3785 VSS.n1491 VSS.n1489 0.237342
R3786 VSS.n1491 VSS.n1490 0.237342
R3787 VSS.n1490 VSS.n318 0.237342
R3788 VSS.n1497 VSS.n318 0.237342
R3789 VSS.n1498 VSS.n1497 0.237342
R3790 VSS.n1501 VSS.n1498 0.237342
R3791 VSS.n1502 VSS.n1501 0.237342
R3792 VSS.n1505 VSS.n1502 0.237342
R3793 VSS.n1506 VSS.n1505 0.237342
R3794 VSS.n1509 VSS.n1506 0.237342
R3795 VSS.n1510 VSS.n1509 0.237342
R3796 VSS.n1515 VSS.n1514 0.237342
R3797 VSS.n1518 VSS.n1515 0.237342
R3798 VSS.n1519 VSS.n1518 0.237342
R3799 VSS.n1520 VSS.n1519 0.237342
R3800 VSS.n1520 VSS.n305 0.237342
R3801 VSS.n1526 VSS.n305 0.237342
R3802 VSS.n1527 VSS.n1526 0.237342
R3803 VSS.n1529 VSS.n1527 0.237342
R3804 VSS.n1529 VSS.n1528 0.237342
R3805 VSS.n1528 VSS.n302 0.237342
R3806 VSS.n1535 VSS.n302 0.237342
R3807 VSS.n1536 VSS.n1535 0.237342
R3808 VSS.n1539 VSS.n1536 0.237342
R3809 VSS.n1540 VSS.n1539 0.237342
R3810 VSS.n1543 VSS.n1540 0.237342
R3811 VSS.n1544 VSS.n1543 0.237342
R3812 VSS.n1547 VSS.n1544 0.237342
R3813 VSS.n1548 VSS.n1547 0.237342
R3814 VSS.n1553 VSS.n1552 0.237342
R3815 VSS.n1556 VSS.n1553 0.237342
R3816 VSS.n1557 VSS.n1556 0.237342
R3817 VSS.n1558 VSS.n1557 0.237342
R3818 VSS.n1558 VSS.n289 0.237342
R3819 VSS.n1564 VSS.n289 0.237342
R3820 VSS.n1565 VSS.n1564 0.237342
R3821 VSS.n1567 VSS.n1565 0.237342
R3822 VSS.n1567 VSS.n1566 0.237342
R3823 VSS.n1566 VSS.n286 0.237342
R3824 VSS.n1574 VSS.n286 0.237342
R3825 VSS.n1575 VSS.n1574 0.237342
R3826 VSS.n1576 VSS.n1575 0.237342
R3827 VSS.n1576 VSS.n284 0.237342
R3828 VSS.n1581 VSS.n284 0.237342
R3829 VSS.n1582 VSS.n1581 0.237342
R3830 VSS.n1582 VSS.n282 0.237342
R3831 VSS.n1587 VSS.n282 0.237342
R3832 VSS.n1634 VSS.n1588 0.237342
R3833 VSS.n1589 VSS.n1588 0.237342
R3834 VSS.n1627 VSS.n1589 0.237342
R3835 VSS.n1627 VSS.n1626 0.237342
R3836 VSS.n1626 VSS.n1625 0.237342
R3837 VSS.n1625 VSS.n1591 0.237342
R3838 VSS.n1620 VSS.n1591 0.237342
R3839 VSS.n1620 VSS.n1619 0.237342
R3840 VSS.n1619 VSS.n1618 0.237342
R3841 VSS.n1618 VSS.n1594 0.237342
R3842 VSS.n1596 VSS.n1594 0.237342
R3843 VSS.n1611 VSS.n1596 0.237342
R3844 VSS.n1611 VSS.n1610 0.237342
R3845 VSS.n1610 VSS.n1609 0.237342
R3846 VSS.n1609 VSS.n1598 0.237342
R3847 VSS.n1604 VSS.n1598 0.237342
R3848 VSS.n1604 VSS.n1603 0.237342
R3849 VSS.n1603 VSS.n1602 0.237342
R3850 VSS.n1900 VSS.n194 0.237342
R3851 VSS.n1900 VSS.n1899 0.237342
R3852 VSS.n1899 VSS.n1898 0.237342
R3853 VSS.n1898 VSS.n197 0.237342
R3854 VSS.n1893 VSS.n197 0.237342
R3855 VSS.n1893 VSS.n1892 0.237342
R3856 VSS.n1892 VSS.n1891 0.237342
R3857 VSS.n1891 VSS.n200 0.237342
R3858 VSS.n204 VSS.n200 0.237342
R3859 VSS.n1885 VSS.n204 0.237342
R3860 VSS.n1885 VSS.n1884 0.237342
R3861 VSS.n1884 VSS.n1883 0.237342
R3862 VSS.n1883 VSS.n205 0.237342
R3863 VSS.n1878 VSS.n205 0.237342
R3864 VSS.n1878 VSS.n1877 0.237342
R3865 VSS.n1877 VSS.n1876 0.237342
R3866 VSS.n1876 VSS.n209 0.237342
R3867 VSS.n1871 VSS.n209 0.237342
R3868 VSS.n1869 VSS.n1856 0.237342
R3869 VSS.n1857 VSS.n1856 0.237342
R3870 VSS.n1862 VSS.n1857 0.237342
R3871 VSS.n1862 VSS.n1861 0.237342
R3872 VSS.n1861 VSS.n1860 0.237342
R3873 VSS.n1860 VSS.n126 0.237342
R3874 VSS.n2031 VSS.n126 0.237342
R3875 VSS.n2032 VSS.n2031 0.237342
R3876 VSS.n2052 VSS.n2032 0.237342
R3877 VSS.n2052 VSS.n2051 0.237342
R3878 VSS.n2051 VSS.n2050 0.237342
R3879 VSS.n2050 VSS.n2033 0.237342
R3880 VSS.n2044 VSS.n2033 0.237342
R3881 VSS.n2044 VSS.n2043 0.237342
R3882 VSS.n2043 VSS.n2042 0.237342
R3883 VSS.n2042 VSS.n2037 0.237342
R3884 VSS.n2037 VSS.n89 0.237342
R3885 VSS.n2188 VSS.n89 0.237342
R3886 VSS.n2191 VSS.n2190 0.237342
R3887 VSS.n2191 VSS.n83 0.237342
R3888 VSS.n2197 VSS.n83 0.237342
R3889 VSS.n2198 VSS.n2197 0.237342
R3890 VSS.n2228 VSS.n2198 0.237342
R3891 VSS.n2228 VSS.n2227 0.237342
R3892 VSS.n2227 VSS.n2226 0.237342
R3893 VSS.n2226 VSS.n2199 0.237342
R3894 VSS.n2220 VSS.n2199 0.237342
R3895 VSS.n2220 VSS.n2219 0.237342
R3896 VSS.n2219 VSS.n2218 0.237342
R3897 VSS.n2218 VSS.n2203 0.237342
R3898 VSS.n2204 VSS.n2203 0.237342
R3899 VSS.n2211 VSS.n2204 0.237342
R3900 VSS.n2211 VSS.n2210 0.237342
R3901 VSS.n2210 VSS.n2209 0.237342
R3902 VSS.n2209 VSS.n23 0.237342
R3903 VSS.n2348 VSS.n23 0.237342
R3904 VSS.n569 VSS.n568 0.237342
R3905 VSS.n569 VSS.n540 0.237342
R3906 VSS.n575 VSS.n540 0.237342
R3907 VSS.n576 VSS.n575 0.237342
R3908 VSS.n577 VSS.n576 0.237342
R3909 VSS.n577 VSS.n536 0.237342
R3910 VSS.n583 VSS.n536 0.237342
R3911 VSS.n584 VSS.n583 0.237342
R3912 VSS.n585 VSS.n584 0.237342
R3913 VSS.n585 VSS.n532 0.237342
R3914 VSS.n591 VSS.n532 0.237342
R3915 VSS.n592 VSS.n591 0.237342
R3916 VSS.n593 VSS.n592 0.237342
R3917 VSS.n593 VSS.n528 0.237342
R3918 VSS.n600 VSS.n528 0.237342
R3919 VSS.n601 VSS.n600 0.237342
R3920 VSS.n2171 VSS.n76 0.237342
R3921 VSS.n2275 VSS.n76 0.237342
R3922 VSS.n2276 VSS.n2275 0.237342
R3923 VSS.n2278 VSS.n2276 0.237342
R3924 VSS.n2278 VSS.n2277 0.237342
R3925 VSS.n2277 VSS.n56 0.237342
R3926 VSS.n695 VSS.n668 0.216026
R3927 VSS.n1222 VSS.n455 0.216026
R3928 VSS.n1390 VSS.n380 0.216026
R3929 VSS.n1303 VSS.n377 0.216026
R3930 VSS.n1434 VSS.n1407 0.216026
R3931 VSS.n1968 VSS.n152 0.216026
R3932 VSS.n1998 VSS.n1997 0.206553
R3933 VSS.n659 VSS.n652 0.192342
R3934 VSS.n1207 VSS.n1206 0.192342
R3935 VSS.n1400 VSS.n383 0.192342
R3936 VSS.n1312 VSS.n378 0.192342
R3937 VSS.n368 VSS.n356 0.192342
R3938 VSS.n1953 VSS.n1952 0.192342
R3939 VSS.n2014 VSS.n141 0.192342
R3940 VSS.n2296 VSS.n55 0.192342
R3941 VSS.n567 VSS.n544 0.192342
R3942 VSS.n111 VSS.n110 0.192342
R3943 VSS.n1163 VSS.n496 0.192342
R3944 VSS.n1770 VSS.n1731 0.192342
R3945 VSS.n249 VSS.n233 0.192342
R3946 VSS.n1036 VSS.n995 0.192342
R3947 VSS.n1071 VSS.n956 0.192342
R3948 VSS.n1106 VSS.n889 0.192342
R3949 VSS.n1206 VSS.n468 0.173395
R3950 VSS.n1400 VSS.n382 0.173395
R3951 VSS.n1269 VSS.n378 0.173395
R3952 VSS.n1281 VSS.n356 0.173395
R3953 VSS.n1952 VSS.n166 0.173395
R3954 VSS.n2014 VSS.n140 0.173395
R3955 VSS.n2296 VSS.n54 0.173395
R3956 VSS.n2298 VSS.n52 0.173395
R3957 VSS.n1163 VSS.n495 0.173395
R3958 VSS.n2072 VSS.n7 0.173395
R3959 VSS.n838 VSS.n835 0.173395
R3960 VSS.n1741 VSS.n1740 0.173395
R3961 VSS.n1726 VSS.n1725 0.173395
R3962 VSS.n1008 VSS.n1007 0.173395
R3963 VSS.n973 VSS.n970 0.173395
R3964 VSS.n906 VSS.n903 0.173395
R3965 VSS.n2173 VSS.n2172 0.161553
R3966 VSS.n603 VSS.n602 0.161553
R3967 VSS.n1157 VSS.n1156 0.161553
R3968 VSS.n1514 VSS.n315 0.161553
R3969 VSS.n1552 VSS.n299 0.161553
R3970 VSS.n1635 VSS.n1634 0.161553
R3971 VSS.n194 VSS.n191 0.161553
R3972 VSS.n1870 VSS.n1869 0.161553
R3973 VSS.n2190 VSS.n2189 0.161553
R3974 VSS.n2316 VSS.n39 0.137868
R3975 VSS VSS.n652 0.124325
R3976 VSS.n2298 VSS.n47 0.119442
R3977 VSS.n703 VSS.n652 0.119442
R3978 VSS.n1158 VSS.n1157 0.114184
R3979 VSS.n1510 VSS.n315 0.114184
R3980 VSS.n1548 VSS.n299 0.114184
R3981 VSS.n1635 VSS.n1587 0.114184
R3982 VSS.n1602 VSS.n191 0.114184
R3983 VSS.n1871 VSS.n1870 0.114184
R3984 VSS.n2189 VSS.n2188 0.114184
R3985 VSS.n2349 VSS.n2348 0.114184
R3986 VSS.n2367 VSS.n2366 0.113
R3987 VSS.n2015 VSS.n2014 0.112898
R3988 VSS.n1952 VSS.n167 0.112898
R3989 VSS.n1442 VSS.n356 0.112898
R3990 VSS.n1375 VSS.n378 0.112898
R3991 VSS.n1400 VSS.n384 0.112898
R3992 VSS.n1206 VSS.n469 0.112898
R3993 VSS.n2296 VSS.n56 0.112898
R3994 VSS.n1222 VSS.n381 0.112876
R3995 VSS.n1404 VSS.n377 0.112876
R3996 VSS.n1968 VSS.n154 0.112876
R3997 VSS.n1407 VSS.n1406 0.112876
R3998 VSS.n1402 VSS.n380 0.112876
R3999 VSS.n668 VSS.n667 0.112876
R4000 VSS.n2189 VSS.n87 0.101158
R4001 VSS.n1870 VSS.n1855 0.101158
R4002 VSS.n1907 VSS.n191 0.101158
R4003 VSS.n1635 VSS.n281 0.101158
R4004 VSS.n1333 VSS.n299 0.101158
R4005 VSS.n404 VSS.n315 0.101158
R4006 VSS.n1157 VSS.n820 0.101158
R4007 VSS.n602 VSS.n526 0.101158
R4008 VSS.n2349 VSS.n22 0.101158
R4009 VSS.n568 VSS.n567 0.100495
R4010 VSS.n2381 VSS.n7 0.100495
R4011 VSS.n2014 VSS.n143 0.0966111
R4012 VSS.n1952 VSS.n169 0.0966111
R4013 VSS.n1405 VSS.n356 0.0966111
R4014 VSS.n1403 VSS.n378 0.0966111
R4015 VSS.n1401 VSS.n1400 0.0966111
R4016 VSS.n1206 VSS.n471 0.0966111
R4017 VSS.n2297 VSS.n2296 0.0966111
R4018 VSS.n1163 VSS.n497 0.0939503
R4019 VSS.n1997 VSS.n53 0.0938027
R4020 VSS.n7 VSS.n1 0.093725
R4021 VSS.n567 VSS 0.089225
R4022 VSS.n2106 VSS.n2105 0.0833947
R4023 VSS.n1777 VSS.n231 0.0833947
R4024 VSS.n1696 VSS.n260 0.0833947
R4025 VSS.n1041 VSS.n994 0.0833947
R4026 VSS.n1076 VSS.n955 0.0833947
R4027 VSS.n1111 VSS.n888 0.0833947
R4028 VSS.n2332 VSS.n2331 0.0798421
R4029 VSS.n2331 VSS.n2330 0.0632632
R4030 VSS.n2189 VSS.n88 0.0466842
R4031 VSS.n1870 VSS.n1810 0.0466842
R4032 VSS.n1662 VSS.n191 0.0466842
R4033 VSS.n1636 VSS.n1635 0.0466842
R4034 VSS.n923 VSS.n299 0.0466842
R4035 VSS.n856 VSS.n315 0.0466842
R4036 VSS.n1157 VSS.n812 0.0466842
R4037 VSS.n2350 VSS.n2349 0.0466842
R4038 VSS.n602 VSS.n601 0.0466842
R4039 VSS.n1163 VSS 0.0446667
R4040 VSS.n689 VSS.n668 0.0443158
R4041 VSS.n1223 VSS.n1222 0.0443158
R4042 VSS.n1384 VSS.n380 0.0443158
R4043 VSS.n1297 VSS.n377 0.0443158
R4044 VSS.n1428 VSS.n1407 0.0443158
R4045 VSS.n1969 VSS.n1968 0.0443158
R4046 VSS.n2368 VSS.n2367 0.0348421
R4047 VSS VSS.n491 0.0307778
R4048 VSS.n143 VSS 0.0307778
R4049 VSS.n169 VSS 0.0307778
R4050 VSS.n1405 VSS 0.0307778
R4051 VSS.n1403 VSS 0.0307778
R4052 VSS.n1401 VSS 0.0307778
R4053 VSS.n471 VSS 0.0307778
R4054 VSS.n2297 VSS 0.0307778
R4055 VSS.n2172 VSS.n2171 0.0289211
R4056 VSS.n2105 VSS 0.0260634
R4057 VSS VSS.n231 0.0260634
R4058 VSS.n260 VSS 0.0260634
R4059 VSS.n1041 VSS 0.0260634
R4060 VSS.n1076 VSS 0.0260634
R4061 VSS.n1111 VSS 0.0260634
R4062 VSS.n2105 VSS.n109 0.0233169
R4063 VSS.n1727 VSS.n231 0.0233169
R4064 VSS.n1006 VSS.n260 0.0233169
R4065 VSS.n1042 VSS.n1041 0.0233169
R4066 VSS.n1077 VSS.n1076 0.0233169
R4067 VSS.n1112 VSS.n1111 0.0233169
R4068 VSS.n1740 VSS.n109 0.0119085
R4069 VSS.n1727 VSS.n1726 0.0119085
R4070 VSS.n1007 VSS.n1006 0.0119085
R4071 VSS.n1042 VSS.n973 0.0119085
R4072 VSS.n1077 VSS.n906 0.0119085
R4073 VSS.n1112 VSS.n838 0.0119085
R4074 VSS.n1997 VSS.n68 0.00997368
R4075 VSS.n2104 VSS.n110 0.00852817
R4076 VSS.n1731 VSS.n1729 0.00852817
R4077 VSS.n259 VSS.n233 0.00852817
R4078 VSS.n1040 VSS.n995 0.00852817
R4079 VSS.n1075 VSS.n956 0.00852817
R4080 VSS.n1110 VSS.n889 0.00852817
R4081 VSS.n2316 VSS.n2315 0.00523684
R4082 VSS VSS.n0 0.00383333
R4083 VSS VSS.n2104 0.0011338
R4084 VSS.n1729 VSS 0.0011338
R4085 VSS VSS.n259 0.0011338
R4086 VSS VSS.n1040 0.0011338
R4087 VSS VSS.n1075 0.0011338
R4088 VSS VSS.n1110 0.0011338
R4089 OUT.n3 OUT.t3 39.434
R4090 OUT.n0 OUT.t5 39.434
R4091 OUT.n3 OUT.t4 29.3205
R4092 OUT.n0 OUT.t2 29.3205
R4093 OUT.n1 OUT.t0 13.7342
R4094 OUT.n2 OUT.n0 8.09525
R4095 OUT.n1 OUT.t1 6.3271
R4096 OUT OUT.n3 1.09775
R4097 OUT.n3 OUT.n2 1.02275
R4098 OUT.n2 OUT.n1 0.3305
R4099 VCNS.n0 VCNS.t3 40.4718
R4100 VCNS.n2 VCNS.t1 40.4081
R4101 VCNS.n1 VCNS.t2 40.4081
R4102 VCNS.n0 VCNS.t0 40.4081
R4103 VCNS VCNS.n2 1.89975
R4104 VCNS.n1 VCNS.n0 0.06425
R4105 VCNS.n2 VCNS.n1 0.06425
R4106 VCNB.n0 VCNB.t2 40.4718
R4107 VCNB.n2 VCNB.t0 40.4081
R4108 VCNB.n1 VCNB.t3 40.4081
R4109 VCNB.n0 VCNB.t1 40.4081
R4110 VCNB VCNB.n2 1.90056
R4111 VCNB.n1 VCNB.n0 0.06425
R4112 VCNB.n2 VCNB.n1 0.06425
R4113 VCTRL VCTRL.t0 29.2551
C0 a_n683_2840 a_n487_2840 0.099479f
C1 a_n8659_n1230 VCNB 0.205658f
C2 a_7177_2840 a_10825_n1138 0.058694f
C3 a_11009_2840 a_10813_2840 0.099479f
C4 a_7177_2840 a_6993_n1138 0.046681f
C5 a_7177_2840 a_10813_2840 0.072091f
C6 a_7177_2840 a_6981_2840 0.099479f
C7 a_7177_2840 a_11009_2840 0.971124f
C8 VDD a_18477_2840 0.298308f
C9 a_18489_n1138 VDD 0.119269f
C10 VDD a_3345_2840 0.629273f
C11 a_14657_n1138 VDD 0.119269f
C12 VDD VCTRL 0.255158f
C13 VDD a_14645_2840 0.298285f
C14 a_10825_n1138 VDD 0.119269f
C15 VDD a_n487_2840 0.629273f
C16 a_6993_n1138 VDD 0.119269f
C17 OUT a_18477_2840 0.073021f
C18 a_18489_n1138 OUT 0.058694f
C19 VDD a_10813_2840 0.298285f
C20 a_3161_n1138 VDD 0.119269f
C21 OUT a_3345_2840 0.142403f
C22 a_14657_n1138 OUT 0.046681f
C23 VDD VCNB 0.307262f
C24 VDD a_6981_2840 0.298285f
C25 a_n671_n1138 VDD 0.119269f
C26 OUT a_14645_2840 0.222712f
C27 a_n8659_n1230 VDD 0.327608f
C28 OUT a_n487_2840 1.12692f
C29 VCTRL a_n9701_6193 0.073173f
C30 VDD a_3149_2840 0.298285f
C31 a_18673_2840 VDD 0.352601f
C32 OUT a_10813_2840 0.122036f
C33 VDD a_n683_2840 0.298285f
C34 a_11009_2840 VDD 0.629273f
C35 OUT a_6981_2840 0.122036f
C36 a_n671_n1138 OUT 0.058694f
C37 a_7177_2840 VDD 0.629273f
C38 OUT a_3149_2840 0.122036f
C39 a_18673_2840 OUT 0.522564f
C40 OUT a_n683_2840 0.198022f
C41 a_11009_2840 OUT 1.11554f
C42 a_7177_2840 OUT 0.142403f
C43 a_n8659_n1230 VCNS 0.1952f
C44 VDD OUT 2.04271f
C45 a_n487_2840 a_3345_2840 0.971124f
C46 a_6993_n1138 a_3345_2840 0.058694f
C47 VDD a_n9701_6193 0.49163f
C48 a_3161_n1138 a_3345_2840 0.046681f
C49 a_6981_2840 a_3345_2840 0.072091f
C50 VDD VCNS 0.35019f
C51 a_18673_2840 a_18477_2840 0.106065f
C52 a_3161_n1138 a_n487_2840 0.058694f
C53 a_18673_2840 a_18489_n1138 0.063905f
C54 a_3149_2840 a_3345_2840 0.099479f
C55 a_n671_n1138 a_n487_2840 0.046681f
C56 a_11009_2840 a_14657_n1138 0.058694f
C57 a_3149_2840 a_n487_2840 0.072091f
C58 a_11009_2840 a_14645_2840 0.072091f
C59 a_7177_2840 a_3345_2840 0.971124f
C60 a_11009_2840 a_10825_n1138 0.046681f
C61 VCNS VSS 2.46604f
C62 VCNB VSS 2.32511f
C63 OUT VSS 13.544005f
C64 VCTRL VSS 2.15234f
C65 VDD VSS 0.133943p
C66 a_18489_n1138 VSS 0.583015f
C67 a_14657_n1138 VSS 0.59026f
C68 a_10825_n1138 VSS 0.59026f
C69 a_6993_n1138 VSS 0.59026f
C70 a_3161_n1138 VSS 0.59026f
C71 a_n671_n1138 VSS 0.59026f
C72 a_n8659_n1230 VSS 2.04692f
C73 a_18673_2840 VSS 1.14559f
C74 a_11009_2840 VSS 3.50221f
C75 a_7177_2840 VSS 3.50221f
C76 a_18477_2840 VSS 0.393424f
C77 a_3345_2840 VSS 3.50221f
C78 a_14645_2840 VSS 0.393424f
C79 a_n487_2840 VSS 3.48363f
C80 a_10813_2840 VSS 0.393424f
C81 a_6981_2840 VSS 0.393424f
C82 a_3149_2840 VSS 0.393424f
C83 a_n683_2840 VSS 0.393424f
C84 a_n9701_6193 VSS 3.02737f
C85 a_16431_6193 VSS 0.776388f
C86 OUT.n0 VSS 0.768913f
C87 OUT.t1 VSS 0.012159f
C88 OUT.n1 VSS 0.077502f
C89 OUT.n2 VSS 0.711343f
C90 OUT.n3 VSS 0.304402f
C91 a_n4208_n141.n0 VSS 0.1651f
C92 a_n4208_n141.n1 VSS 2.04471f
C93 a_n4208_n141.n2 VSS 0.898532f
C94 a_n4208_n141.n3 VSS 1.1521f
C95 a_n4208_n141.t4 VSS 0.026172f
C96 a_n4208_n141.t2 VSS 0.068133f
C97 VDD.t17 VSS 0.056965f
C98 VDD.n2 VSS 0.038057f
C99 VDD.t21 VSS 0.079048f
C100 VDD.n3 VSS 0.078931f
C101 VDD.n5 VSS 0.106518f
C102 VDD.t9 VSS 0.056965f
C103 VDD.n8 VSS 0.038057f
C104 VDD.t0 VSS 0.079048f
C105 VDD.n9 VSS 0.078931f
C106 VDD.n11 VSS 0.056372f
C107 VDD.n12 VSS 0.182172f
C108 VDD.t5 VSS 0.056965f
C109 VDD.n15 VSS 0.038057f
C110 VDD.t3 VSS 0.079048f
C111 VDD.n16 VSS 0.078931f
C112 VDD.n18 VSS 0.056372f
C113 VDD.n19 VSS 0.181181f
C114 VDD.t7 VSS 0.056965f
C115 VDD.n22 VSS 0.038057f
C116 VDD.t4 VSS 0.079048f
C117 VDD.n23 VSS 0.078931f
C118 VDD.n25 VSS 0.056372f
C119 VDD.n26 VSS 0.181181f
C120 VDD.t19 VSS 0.056965f
C121 VDD.n29 VSS 0.038057f
C122 VDD.t2 VSS 0.079048f
C123 VDD.n30 VSS 0.078931f
C124 VDD.n32 VSS 0.056372f
C125 VDD.n33 VSS 0.181181f
C126 VDD.t13 VSS 0.056965f
C127 VDD.n36 VSS 0.038057f
C128 VDD.t1 VSS 0.079048f
C129 VDD.n37 VSS 0.078931f
C130 VDD.n39 VSS 0.056372f
C131 VDD.n40 VSS 0.181181f
C132 VDD.t11 VSS 0.056965f
C133 VDD.n41 VSS 0.060525f
C134 VDD.t15 VSS 0.056965f
C135 VDD.n42 VSS 0.063689f
C136 VDD.n43 VSS 0.092744f
C137 VDD.n44 VSS 0.232621f
C138 a_n8471_219.n0 VSS 3.08842f
C139 a_n8471_219.n1 VSS 1.16302f
C140 a_n8471_219.n2 VSS 1.4992f
C141 a_n8471_219.n3 VSS 0.343638f
C142 a_n8471_219.t2 VSS 0.038537f
C143 a_n8471_219.t1 VSS 0.039863f
C144 a_n8471_219.t4 VSS 0.013068f
C145 a_n8471_219.t8 VSS 0.01284f
C146 a_n8471_219.t6 VSS 0.031089f
C147 a_n8471_219.t9 VSS 0.011094f
C148 a_n8471_219.t11 VSS 0.011094f
C149 a_n8471_219.t10 VSS 0.011094f
C150 a_n8471_219.t5 VSS 0.011094f
C151 a_n8471_219.t7 VSS 0.011094f
C152 a_n8471_219.t0 VSS 0.024053f
C153 a_n8471_219.n4 VSS 0.382885f
.ends

