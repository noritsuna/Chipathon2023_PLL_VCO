* NGSPICE file created from TOP.ext - technology: gf180mcuD

.subckt TOP VDD OUT vctrl VCNB VCNS VSS
X0 VSS a_n4208_n113# a_n671_n1136# VSS nfet_03v3 ad=0.427p pd=2.62u as=0.427p ps=2.62u w=0.7u l=0.33u
X1 VDD a_n8471_219# a_3149_2840# VDD pfet_03v3 ad=1.17p pd=4.9u as=1.17p ps=4.9u w=1.8u l=0.33u
X2 a_7177_2840# a_3345_2840# a_6981_2840# VDD pfet_03v3 ad=2.34p pd=8.5u as=2.34p ps=8.5u w=3.6u l=0.33u
X3 VSS VCNS a_n8659_n1230# VSS nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.33u
X4 a_n9701_6793# a_16431_6193# VSS ppolyf_u r_width=0.8u r_length=0.13m
X5 a_n8471_219# VCNB a_n8659_n1230# VSS nfet_03v3 ad=0.52p pd=2.52u as=1.22p ps=5.22u w=2u l=0.33u
X6 VDD a_n8471_219# a_n8471_219# VDD pfet_03v3 ad=1.17p pd=4.9u as=1.17p ps=4.9u w=1.8u l=0.33u
X7 VDD a_n8471_219# a_18477_2840# VDD pfet_03v3 ad=1.17p pd=4.9u as=1.17p ps=4.9u w=1.8u l=0.33u
X8 VSS VCNS a_n8659_n1230# VSS nfet_03v3 ad=0.52p pd=2.52u as=1.22p ps=5.22u w=2u l=0.33u
X9 VDD a_n8471_219# a_n683_2840# VDD pfet_03v3 ad=1.17p pd=4.9u as=1.17p ps=4.9u w=1.8u l=0.33u
X10 a_11009_2840# a_7177_2840# a_10813_2840# VDD pfet_03v3 ad=2.34p pd=8.5u as=2.34p ps=8.5u w=3.6u l=0.33u
X11 a_n487_2840# OUT a_n671_n1136# VSS nfet_03v3 ad=0.854p pd=4.02u as=0.854p ps=4.02u w=1.4u l=0.33u
X12 a_7177_2840# a_3345_2840# a_6993_n1136# VSS nfet_03v3 ad=0.854p pd=4.02u as=0.854p ps=4.02u w=1.4u l=0.33u
X13 a_n9701_6793# a_16431_7393# VSS ppolyf_u r_width=0.8u r_length=0.13m
X14 a_3345_2840# a_n487_2840# a_3149_2840# VDD pfet_03v3 ad=2.34p pd=8.5u as=2.34p ps=8.5u w=3.6u l=0.33u
X15 a_18673_2840# OUT a_18489_n1136# VSS nfet_03v3 ad=0.854p pd=4.02u as=0.854p ps=4.02u w=1.4u l=0.33u
X16 VSS a_16431_7393# VSS ppolyf_u r_width=0.8u r_length=0.13m
X17 a_n8471_219# vctrl a_n9701_6193# VSS nfet_03v3 ad=0.488p pd=2.82u as=0.488p ps=2.82u w=0.8u l=0.33u
X18 a_18673_2840# OUT a_18477_2840# VDD pfet_03v3 ad=2.34p pd=8.5u as=2.34p ps=8.5u w=3.6u l=0.33u
X19 VSS a_n4208_n113# a_18489_n1136# VSS nfet_03v3 ad=0.427p pd=2.62u as=0.427p ps=2.62u w=0.7u l=0.33u
X20 a_n487_2840# OUT a_n683_2840# VDD pfet_03v3 ad=2.34p pd=8.5u as=2.34p ps=8.5u w=3.6u l=0.33u
X21 a_n8659_n1230# VCNS VSS VSS nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.33u
X22 VDD a_n8471_219# a_14645_2840# VDD pfet_03v3 ad=1.17p pd=4.9u as=1.17p ps=4.9u w=1.8u l=0.33u
X23 VSS a_n4208_n113# a_14657_n1136# VSS nfet_03v3 ad=0.427p pd=2.62u as=0.427p ps=2.62u w=0.7u l=0.33u
X24 a_n4208_n113# a_n8471_219# VDD VDD pfet_03v3 ad=1.17p pd=4.9u as=1.17p ps=4.9u w=1.8u l=0.33u
X25 a_11009_2840# a_7177_2840# a_10825_n1136# VSS nfet_03v3 ad=0.854p pd=4.02u as=0.854p ps=4.02u w=1.4u l=0.33u
X26 VSS a_n4208_n113# a_3161_n1136# VSS nfet_03v3 ad=0.427p pd=2.62u as=0.427p ps=2.62u w=0.7u l=0.33u
X27 a_n8471_219# VCNB a_n8659_n1230# VSS nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.33u
X28 VDD a_n8471_219# a_6981_2840# VDD pfet_03v3 ad=1.17p pd=4.9u as=1.17p ps=4.9u w=1.8u l=0.33u
X29 a_3345_2840# a_n487_2840# a_3161_n1136# VSS nfet_03v3 ad=0.854p pd=4.02u as=0.854p ps=4.02u w=1.4u l=0.33u
X30 VSS a_n4208_n113# a_6993_n1136# VSS nfet_03v3 ad=0.427p pd=2.62u as=0.427p ps=2.62u w=0.7u l=0.33u
X31 a_n8659_n1230# VCNB a_n8471_219# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.52p ps=2.52u w=2u l=0.33u
X32 a_n8659_n1230# VCNS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0.52p ps=2.52u w=2u l=0.33u
X33 VSS a_n4208_n113# a_10825_n1136# VSS nfet_03v3 ad=0.427p pd=2.62u as=0.427p ps=2.62u w=0.7u l=0.33u
X34 a_n4208_n113# a_n4208_n113# VSS VSS nfet_03v3 ad=0.427p pd=2.62u as=0.427p ps=2.62u w=0.7u l=0.33u
X35 a_n9701_6193# a_16431_6193# VSS ppolyf_u r_width=0.8u r_length=0.13m
X36 a_n8659_n1230# VCNB a_n8471_219# VSS nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.33u
X37 OUT a_11009_2840# a_14657_n1136# VSS nfet_03v3 ad=0.854p pd=4.02u as=0.854p ps=4.02u w=1.4u l=0.33u
X38 VDD a_n8471_219# a_10813_2840# VDD pfet_03v3 ad=1.17p pd=4.9u as=1.17p ps=4.9u w=1.8u l=0.33u
X39 OUT a_11009_2840# a_14645_2840# VDD pfet_03v3 ad=2.34p pd=8.5u as=2.34p ps=8.5u w=3.6u l=0.33u
C0 a_n8659_n1230# VCNS 0.1952f
C1 a_n487_2840# VDD 0.790856f
C2 VDD a_n8471_219# 6.43873f
C3 a_18477_2840# a_n8471_219# 0.034056f
C4 a_n9701_6193# a_n8471_219# 0.030193f
C5 a_n487_2840# a_n683_2840# 0.239058f
C6 a_n671_n1136# OUT 0.063619f
C7 a_n8471_219# a_n683_2840# 0.032842f
C8 a_18489_n1136# OUT 0.063703f
C9 a_18673_2840# a_n8471_219# 8.34e-20
C10 a_3149_2840# a_3345_2840# 0.239058f
C11 a_3345_2840# a_n4208_n113# 8.03e-19
C12 a_6981_2840# a_3345_2840# 0.105347f
C13 a_3149_2840# OUT 0.126347f
C14 a_18477_2840# VDD 0.297366f
C15 OUT a_n4208_n113# 0.108655f
C16 a_6993_n1136# a_7177_2840# 0.067104f
C17 a_10825_n1136# a_n4208_n113# 0.013607f
C18 a_6981_2840# OUT 0.126347f
C19 a_11009_2840# a_n4208_n113# 8.03e-19
C20 a_16431_6193# a_n8471_219# 2.66e-19
C21 a_n9701_6193# VDD 0.406316f
C22 VDD a_n683_2840# 0.297325f
C23 a_n487_2840# a_3161_n1136# 0.063619f
C24 a_18673_2840# VDD 0.633399f
C25 a_18477_2840# a_18673_2840# 0.253072f
C26 VCNB a_n8471_219# 0.194241f
C27 a_n487_2840# a_n671_n1136# 0.067104f
C28 a_16431_6193# VDD 0.0038f
C29 a_7177_2840# a_n4208_n113# 8.03e-19
C30 a_3345_2840# OUT 0.161349f
C31 a_6981_2840# a_7177_2840# 0.239058f
C32 a_3149_2840# a_n487_2840# 0.105347f
C33 VCNB VDD 0.115897f
C34 a_14645_2840# OUT 0.365796f
C35 a_3149_2840# a_n8471_219# 0.032842f
C36 a_n487_2840# a_n4208_n113# 8.03e-19
C37 a_n8471_219# a_n4208_n113# 0.034668f
C38 a_11009_2840# OUT 1.09417f
C39 a_10825_n1136# a_11009_2840# 0.067104f
C40 a_11009_2840# a_14645_2840# 0.105347f
C41 a_n8659_n1230# a_n8471_219# 0.691294f
C42 a_14657_n1136# a_n4208_n113# 0.013607f
C43 a_6981_2840# a_n8471_219# 0.032842f
C44 VCNS a_n8471_219# 0.001233f
C45 a_16431_6193# a_16431_7393# 0.010032f
C46 a_18489_n1136# a_18673_2840# 0.071243f
C47 a_3345_2840# a_7177_2840# 0.930892f
C48 a_3149_2840# VDD 0.297325f
C49 VDD a_n4208_n113# 3.44655f
C50 a_10813_2840# OUT 0.126347f
C51 a_n8659_n1230# VDD 7.43e-19
C52 a_6981_2840# VDD 0.297325f
C53 a_10813_2840# a_11009_2840# 0.239058f
C54 OUT a_7177_2840# 0.161349f
C55 a_10825_n1136# a_7177_2840# 0.063619f
C56 a_n487_2840# a_3345_2840# 0.930892f
C57 a_11009_2840# a_7177_2840# 0.930892f
C58 a_3345_2840# a_n8471_219# 0.002936f
C59 VCNS VDD 0.199523f
C60 a_18673_2840# a_n4208_n113# 9.22e-21
C61 a_n487_2840# OUT 1.119f
C62 a_n8471_219# OUT 0.873835f
C63 a_n8471_219# a_14645_2840# 0.032842f
C64 a_14657_n1136# OUT 0.067104f
C65 a_11009_2840# a_n8471_219# 0.002936f
C66 a_14657_n1136# a_11009_2840# 0.063619f
C67 a_n9701_6193# a_n9701_6793# 0.015999f
C68 VDD a_3345_2840# 0.790856f
C69 a_10813_2840# a_7177_2840# 0.105347f
C70 a_3161_n1136# a_n4208_n113# 0.013607f
C71 a_6993_n1136# a_n4208_n113# 0.013607f
C72 VDD OUT 2.27325f
C73 a_18477_2840# OUT 0.106543f
C74 VDD a_14645_2840# 0.297325f
C75 a_11009_2840# VDD 0.790856f
C76 a_10813_2840# a_n8471_219# 0.032842f
C77 a_n8659_n1230# VCNB 0.205658f
C78 a_n8471_219# vctrl 0.007799f
C79 a_n8471_219# a_7177_2840# 0.002936f
C80 a_n683_2840# OUT 0.236339f
C81 a_n671_n1136# a_n4208_n113# 0.013607f
C82 a_18673_2840# OUT 0.566131f
C83 VCNB VCNS 0.003188f
C84 a_18489_n1136# a_n4208_n113# 0.013607f
C85 a_n487_2840# a_n8471_219# 0.002936f
C86 a_3345_2840# a_3161_n1136# 0.067104f
C87 a_10813_2840# VDD 0.297325f
C88 VDD vctrl 0.130527f
C89 a_3345_2840# a_6993_n1136# 0.063619f
C90 VDD a_7177_2840# 0.790856f
C91 a_n9701_6193# vctrl 0.073173f
C92 VCNS VSS 2.63992f
C93 VCNB VSS 2.51968f
C94 OUT VSS 13.4135f
C95 vctrl VSS 2.27922f
C96 VDD VSS 81.2828f
C97 a_18489_n1136# VSS 0.747362f
C98 a_14657_n1136# VSS 0.747362f
C99 a_10825_n1136# VSS 0.747362f
C100 a_6993_n1136# VSS 0.747362f
C101 a_3161_n1136# VSS 0.747362f
C102 a_n671_n1136# VSS 0.747362f
C103 a_n8659_n1230# VSS 2.37379f
C104 a_18673_2840# VSS 1.32356f
C105 a_11009_2840# VSS 3.71444f
C106 a_18477_2840# VSS 0.292039f
C107 a_7177_2840# VSS 3.71444f
C108 a_14645_2840# VSS 0.292039f
C109 a_3345_2840# VSS 3.71444f
C110 a_10813_2840# VSS 0.292039f
C111 a_n487_2840# VSS 3.67709f
C112 a_6981_2840# VSS 0.292039f
C113 a_3149_2840# VSS 0.292039f
C114 a_n4208_n113# VSS 21.5682f
C115 a_n683_2840# VSS 0.292039f
C116 a_n8471_219# VSS 15.745701f
C117 a_n9701_6193# VSS 3.09512f
C118 a_16431_6193# VSS 0.768771f
C119 a_n9701_6793# VSS 0.835507f
C120 a_16431_7393# VSS 0.76357f
.ends

