* Extracted by KLayout with GF180MCU LVS runset on : 09/01/2024 13:11

.SUBCKT TOP VSS VCTRL OUT VCNB VCNS
R$1 \$8 VSS VSS 113750 ppolyf_u L=260U W=0.8U
M$3 VSS VCNS \$7 VSS nfet_03v3_dn L=0.33U W=8U AS=2.78P AD=2.78P PS=12.78U
+ PD=12.78U
M$7 \$10 VCNB \$7 VSS nfet_03v3_dn L=0.33U W=8U AS=2.78P AD=2.78P PS=12.78U
+ PD=12.78U
M$11 \$8 VCTRL \$10 VSS nfet_03v3_dn L=0.33U W=0.8U AS=0.488P AD=0.488P
+ PS=2.82U PD=2.82U
M$12 \$6 \$10 \$11 \$6 pfet_03v3 L=0.33U W=0.9U AS=0.585P AD=0.585P PS=3.1U
+ PD=3.1U
M$13 VSS \$11 \$11 VSS nfet_03v3_dn L=0.33U W=0.42U AS=0.2646P AD=0.2646P
+ PS=2.1U PD=2.1U
M$14 VSS \$11 \$I142 VSS nfet_03v3_dn L=0.33U W=0.42U AS=0.2646P AD=0.2646P
+ PS=2.1U PD=2.1U
M$15 VSS \$11 \$I154 VSS nfet_03v3_dn L=0.33U W=0.42U AS=0.2646P AD=0.2646P
+ PS=2.1U PD=2.1U
M$16 VSS \$11 \$I167 VSS nfet_03v3_dn L=0.33U W=0.42U AS=0.2646P AD=0.2646P
+ PS=2.1U PD=2.1U
M$17 VSS \$11 \$I180 VSS nfet_03v3_dn L=0.33U W=0.42U AS=0.2646P AD=0.2646P
+ PS=2.1U PD=2.1U
M$18 VSS \$11 \$I193 VSS nfet_03v3_dn L=0.33U W=0.42U AS=0.2646P AD=0.2646P
+ PS=2.1U PD=2.1U
M$19 VSS \$11 \$I206 VSS nfet_03v3_dn L=0.33U W=0.42U AS=0.2646P AD=0.2646P
+ PS=2.1U PD=2.1U
M$20 \$I140 OUT \$I146 \$6 pfet_03v3 L=0.33U W=1.8U AS=1.17P AD=1.17P PS=4.9U
+ PD=4.9U
M$21 \$I63 \$I71 \$I159 \$6 pfet_03v3 L=0.33U W=1.8U AS=1.17P AD=1.17P PS=4.9U
+ PD=4.9U
M$22 \$I71 OUT \$I172 \$6 pfet_03v3 L=0.33U W=1.8U AS=1.17P AD=1.17P PS=4.9U
+ PD=4.9U
M$23 \$I64 \$I63 \$I185 \$6 pfet_03v3 L=0.33U W=1.8U AS=1.17P AD=1.17P PS=4.9U
+ PD=4.9U
M$24 \$I65 \$I64 \$I198 \$6 pfet_03v3 L=0.33U W=1.8U AS=1.17P AD=1.17P PS=4.9U
+ PD=4.9U
M$25 OUT \$I65 \$I211 \$6 pfet_03v3 L=0.33U W=1.8U AS=1.17P AD=1.17P PS=4.9U
+ PD=4.9U
M$26 \$6 \$10 \$10 \$6 pfet_03v3 L=0.33U W=0.9U AS=0.585P AD=0.585P PS=3.1U
+ PD=3.1U
M$27 \$6 \$10 \$I146 \$6 pfet_03v3 L=0.33U W=0.9U AS=0.585P AD=0.585P PS=3.1U
+ PD=3.1U
M$28 \$6 \$10 \$I159 \$6 pfet_03v3 L=0.33U W=0.9U AS=0.585P AD=0.585P PS=3.1U
+ PD=3.1U
M$29 \$6 \$10 \$I172 \$6 pfet_03v3 L=0.33U W=0.9U AS=0.585P AD=0.585P PS=3.1U
+ PD=3.1U
M$30 \$6 \$10 \$I185 \$6 pfet_03v3 L=0.33U W=0.9U AS=0.585P AD=0.585P PS=3.1U
+ PD=3.1U
M$31 \$6 \$10 \$I198 \$6 pfet_03v3 L=0.33U W=0.9U AS=0.585P AD=0.585P PS=3.1U
+ PD=3.1U
M$32 \$6 \$10 \$I211 \$6 pfet_03v3 L=0.33U W=0.9U AS=0.585P AD=0.585P PS=3.1U
+ PD=3.1U
M$33 \$I140 OUT \$I142 VSS nfet_03v3_dn L=0.33U W=0.84U AS=0.5124P AD=0.5124P
+ PS=2.9U PD=2.9U
M$34 \$I63 \$I71 \$I154 VSS nfet_03v3_dn L=0.33U W=0.84U AS=0.5124P AD=0.5124P
+ PS=2.9U PD=2.9U
M$35 \$I71 OUT \$I167 VSS nfet_03v3_dn L=0.33U W=0.84U AS=0.5124P AD=0.5124P
+ PS=2.9U PD=2.9U
M$36 \$I64 \$I63 \$I180 VSS nfet_03v3_dn L=0.33U W=0.84U AS=0.5124P AD=0.5124P
+ PS=2.9U PD=2.9U
M$37 \$I65 \$I64 \$I193 VSS nfet_03v3_dn L=0.33U W=0.84U AS=0.5124P AD=0.5124P
+ PS=2.9U PD=2.9U
M$38 OUT \$I65 \$I206 VSS nfet_03v3_dn L=0.33U W=0.84U AS=0.5124P AD=0.5124P
+ PS=2.9U PD=2.9U
.ENDS TOP
