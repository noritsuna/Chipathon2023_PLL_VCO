* NGSPICE file created from TOP.ext - technology: gf180mcuD

.subckt TOP VDD OUT vctrl VCNB VCNS VSS
X0 VSS a_n4208_n113 a_n671_n1136 VSS nfet_03v3 ad=0.427p pd=2.62u as=0.427p ps=2.62u w=0.7u l=0.33u
X1 VDD a_n8471_219 a_3149_2840 VDD pfet_03v3 ad=1.17p pd=4.9u as=1.17p ps=4.9u w=1.8u l=0.33u
X2 a_7177_2840 a_3345_2840 a_6981_2840 VDD pfet_03v3 ad=2.34p pd=8.5u as=2.34p ps=8.5u w=3.6u l=0.33u
X3 VSS VCNS a_n8659_n1230 VSS nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.33u
X4 a_n9701_6793 a_16431_6193 VSS ppolyf_u r_width=0.8u r_length=0.13m
X5 a_n8471_219 VCNB a_n8659_n1230 VSS nfet_03v3 ad=0.52p pd=2.52u as=1.22p ps=5.22u w=2u l=0.33u
X6 VDD a_n8471_219 a_n8471_219 VDD pfet_03v3 ad=1.17p pd=4.9u as=1.17p ps=4.9u w=1.8u l=0.33u
X7 VDD a_n8471_219 a_18477_2840 VDD pfet_03v3 ad=1.17p pd=4.9u as=1.17p ps=4.9u w=1.8u l=0.33u
X8 VSS VCNS a_n8659_n1230 VSS nfet_03v3 ad=0.52p pd=2.52u as=1.22p ps=5.22u w=2u l=0.33u
X9 VDD a_n8471_219 a_n683_2840 VDD pfet_03v3 ad=1.17p pd=4.9u as=1.17p ps=4.9u w=1.8u l=0.33u
X10 a_11009_2840 a_7177_2840 a_10813_2840 VDD pfet_03v3 ad=2.34p pd=8.5u as=2.34p ps=8.5u w=3.6u l=0.33u
X11 a_n487_2840 OUT a_n671_n1136 VSS nfet_03v3 ad=0.854p pd=4.02u as=0.854p ps=4.02u w=1.4u l=0.33u
X12 a_7177_2840 a_3345_2840 a_6993_n1136 VSS nfet_03v3 ad=0.854p pd=4.02u as=0.854p ps=4.02u w=1.4u l=0.33u
X13 a_n9701_6793 a_16431_7393 VSS ppolyf_u r_width=0.8u r_length=0.13m
X14 a_3345_2840 a_n487_2840 a_3149_2840 VDD pfet_03v3 ad=2.34p pd=8.5u as=2.34p ps=8.5u w=3.6u l=0.33u
X15 a_18673_2840 OUT a_18489_n1136 VSS nfet_03v3 ad=0.854p pd=4.02u as=0.854p ps=4.02u w=1.4u l=0.33u
X16 VSS a_16431_7393 VSS ppolyf_u r_width=0.8u r_length=0.13m
X17 a_n8471_219 vctrl a_n9701_6193 VSS nfet_03v3 ad=0.488p pd=2.82u as=0.488p ps=2.82u w=0.8u l=0.33u
X18 a_18673_2840 OUT a_18477_2840 VDD pfet_03v3 ad=2.34p pd=8.5u as=2.34p ps=8.5u w=3.6u l=0.33u
X19 VSS a_n4208_n113 a_18489_n1136 VSS nfet_03v3 ad=0.427p pd=2.62u as=0.427p ps=2.62u w=0.7u l=0.33u
X20 a_n487_2840 OUT a_n683_2840 VDD pfet_03v3 ad=2.34p pd=8.5u as=2.34p ps=8.5u w=3.6u l=0.33u
X21 a_n8659_n1230 VCNS VSS VSS nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.33u
X22 VDD a_n8471_219 a_14645_2840 VDD pfet_03v3 ad=1.17p pd=4.9u as=1.17p ps=4.9u w=1.8u l=0.33u
X23 VSS a_n4208_n113 a_14657_n1136 VSS nfet_03v3 ad=0.427p pd=2.62u as=0.427p ps=2.62u w=0.7u l=0.33u
X24 a_n4208_n113 a_n8471_219 VDD VDD pfet_03v3 ad=1.17p pd=4.9u as=1.17p ps=4.9u w=1.8u l=0.33u
X25 a_11009_2840 a_7177_2840 a_10825_n1136 VSS nfet_03v3 ad=0.854p pd=4.02u as=0.854p ps=4.02u w=1.4u l=0.33u
X26 VSS a_n4208_n113 a_3161_n1136 VSS nfet_03v3 ad=0.427p pd=2.62u as=0.427p ps=2.62u w=0.7u l=0.33u
X27 a_n8471_219 VCNB a_n8659_n1230 VSS nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.33u
X28 VDD a_n8471_219 a_6981_2840 VDD pfet_03v3 ad=1.17p pd=4.9u as=1.17p ps=4.9u w=1.8u l=0.33u
X29 a_3345_2840 a_n487_2840 a_3161_n1136 VSS nfet_03v3 ad=0.854p pd=4.02u as=0.854p ps=4.02u w=1.4u l=0.33u
X30 VSS a_n4208_n113 a_6993_n1136 VSS nfet_03v3 ad=0.427p pd=2.62u as=0.427p ps=2.62u w=0.7u l=0.33u
X31 a_n8659_n1230 VCNB a_n8471_219 VSS nfet_03v3 ad=1.22p pd=5.22u as=0.52p ps=2.52u w=2u l=0.33u
X32 a_n8659_n1230 VCNS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0.52p ps=2.52u w=2u l=0.33u
X33 VSS a_n4208_n113 a_10825_n1136 VSS nfet_03v3 ad=0.427p pd=2.62u as=0.427p ps=2.62u w=0.7u l=0.33u
X34 a_n4208_n113 a_n4208_n113 VSS VSS nfet_03v3 ad=0.427p pd=2.62u as=0.427p ps=2.62u w=0.7u l=0.33u
X35 a_n9701_6193 a_16431_6193 VSS ppolyf_u r_width=0.8u r_length=0.13m
X36 a_n8659_n1230 VCNB a_n8471_219 VSS nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.33u
X37 OUT a_11009_2840 a_14657_n1136 VSS nfet_03v3 ad=0.854p pd=4.02u as=0.854p ps=4.02u w=1.4u l=0.33u
X38 VDD a_n8471_219 a_10813_2840 VDD pfet_03v3 ad=1.17p pd=4.9u as=1.17p ps=4.9u w=1.8u l=0.33u
X39 OUT a_11009_2840 a_14645_2840 VDD pfet_03v3 ad=2.34p pd=8.5u as=2.34p ps=8.5u w=3.6u l=0.33u
C0 a_n4208_n113 a_n8471_219 0.034668f
C1 VDD a_n4208_n113 3.44655f
C2 a_11009_2840 a_n4208_n113 8.03e-19
C3 OUT a_n671_n1136 0.063619f
C4 OUT a_6981_2840 0.126347f
C5 a_n8659_n1230 a_n8471_219 0.691294f
C6 a_3345_2840 a_3161_n1136 0.067104f
C7 VDD a_n8659_n1230 7.43e-19
C8 a_18489_n1136 a_n4208_n113 0.013607f
C9 a_18673_2840 a_n8471_219 8.34e-20
C10 a_n4208_n113 a_3345_2840 8.03e-19
C11 VDD a_18673_2840 0.633399f
C12 a_n4208_n113 a_14657_n1136 0.013607f
C13 VCNB a_n8471_219 0.194241f
C14 VDD VCNB 0.115897f
C15 a_18489_n1136 a_18673_2840 0.071243f
C16 a_n4208_n113 a_3161_n1136 0.013607f
C17 a_7177_2840 a_n8471_219 0.002936f
C18 VDD a_7177_2840 0.790856f
C19 a_3345_2840 a_6993_n1136 0.063619f
C20 a_n487_2840 a_n8471_219 0.002936f
C21 a_11009_2840 a_7177_2840 0.930892f
C22 VCNS a_n8659_n1230 0.1952f
C23 VDD a_n487_2840 0.790856f
C24 a_3149_2840 a_n487_2840 0.105347f
C25 a_7177_2840 a_3345_2840 0.930892f
C26 OUT a_n8471_219 0.873835f
C27 VDD OUT 2.27325f
C28 a_n4208_n113 a_18673_2840 9.22e-21
C29 a_n487_2840 a_3345_2840 0.930892f
C30 VCNS VCNB 0.003188f
C31 OUT a_11009_2840 1.09417f
C32 a_n4208_n113 a_6993_n1136 0.013607f
C33 OUT a_3149_2840 0.126347f
C34 a_18489_n1136 OUT 0.063703f
C35 OUT a_3345_2840 0.161349f
C36 OUT a_14657_n1136 0.067104f
C37 a_n487_2840 a_3161_n1136 0.063619f
C38 a_n4208_n113 a_7177_2840 8.03e-19
C39 VCNB a_n8659_n1230 0.205658f
C40 vctrl a_n9701_6193 0.073173f
C41 vctrl a_n8471_219 0.007799f
C42 a_n487_2840 a_n4208_n113 8.03e-19
C43 a_16431_7393 a_16431_6193 0.010032f
C44 VDD vctrl 0.130527f
C45 a_14645_2840 a_n8471_219 0.032842f
C46 VDD a_14645_2840 0.297325f
C47 a_11009_2840 a_14645_2840 0.105347f
C48 a_10813_2840 a_n8471_219 0.032842f
C49 OUT a_n4208_n113 0.108655f
C50 a_n683_2840 a_n8471_219 0.032842f
C51 VDD a_10813_2840 0.297325f
C52 VDD a_n683_2840 0.297325f
C53 a_7177_2840 a_6993_n1136 0.067104f
C54 a_10813_2840 a_11009_2840 0.239058f
C55 a_18477_2840 a_n8471_219 0.034056f
C56 VDD a_18477_2840 0.297366f
C57 OUT a_18673_2840 0.566131f
C58 OUT a_7177_2840 0.161349f
C59 a_6981_2840 a_n8471_219 0.032842f
C60 OUT a_n487_2840 1.119f
C61 a_11009_2840 a_10825_n1136 0.067104f
C62 VDD a_6981_2840 0.297325f
C63 a_6981_2840 a_3345_2840 0.105347f
C64 a_16431_6193 a_n8471_219 2.66e-19
C65 a_18477_2840 a_18673_2840 0.253072f
C66 VDD a_16431_6193 0.0038f
C67 a_10813_2840 a_7177_2840 0.105347f
C68 a_n4208_n113 a_10825_n1136 0.013607f
C69 a_n4208_n113 a_n671_n1136 0.013607f
C70 a_n683_2840 a_n487_2840 0.239058f
C71 a_n9701_6193 a_n8471_219 0.030193f
C72 VDD a_n9701_6193 0.406316f
C73 OUT a_14645_2840 0.365796f
C74 VDD a_n8471_219 6.43873f
C75 a_11009_2840 a_n8471_219 0.002936f
C76 OUT a_10813_2840 0.126347f
C77 OUT a_n683_2840 0.236339f
C78 VDD a_11009_2840 0.790856f
C79 a_3149_2840 a_n8471_219 0.032842f
C80 VDD a_3149_2840 0.297325f
C81 a_3345_2840 a_n8471_219 0.002936f
C82 VDD a_3345_2840 0.790856f
C83 OUT a_18477_2840 0.106543f
C84 a_7177_2840 a_10825_n1136 0.063619f
C85 a_11009_2840 a_14657_n1136 0.063619f
C86 a_3149_2840 a_3345_2840 0.239058f
C87 a_6981_2840 a_7177_2840 0.239058f
C88 VCNS a_n8471_219 0.001233f
C89 VDD VCNS 0.199523f
C90 a_n487_2840 a_n671_n1136 0.067104f
C91 a_n9701_6793 a_n9701_6193 0.015999f
C92 VCNS VSS 2.63992f
C93 VCNB VSS 2.51968f
C94 OUT VSS 13.4135f
C95 vctrl VSS 2.27922f
C96 VDD VSS 81.2828f
C97 a_18489_n1136 VSS 0.747362f
C98 a_14657_n1136 VSS 0.747362f
C99 a_10825_n1136 VSS 0.747362f
C100 a_6993_n1136 VSS 0.747362f
C101 a_3161_n1136 VSS 0.747362f
C102 a_n671_n1136 VSS 0.747362f
C103 a_n8659_n1230 VSS 2.37379f
C104 a_18673_2840 VSS 1.32356f
C105 a_11009_2840 VSS 3.71444f
C106 a_18477_2840 VSS 0.292039f
C107 a_7177_2840 VSS 3.71444f
C108 a_14645_2840 VSS 0.292039f
C109 a_3345_2840 VSS 3.71444f
C110 a_10813_2840 VSS 0.292039f
C111 a_n487_2840 VSS 3.67709f
C112 a_6981_2840 VSS 0.292039f
C113 a_3149_2840 VSS 0.292039f
C114 a_n4208_n113 VSS 21.5682f
C115 a_n683_2840 VSS 0.292039f
C116 a_n8471_219 VSS 15.745701f
C117 a_n9701_6193 VSS 3.09512f
C118 a_16431_6193 VSS 0.768771f
C119 a_n9701_6793 VSS 0.835507f
C120 a_16431_7393 VSS 0.76357f
.ends

